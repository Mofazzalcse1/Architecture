CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
210 400 30 70 10
176 80 1364 699
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
177
13 Logic Switch~
5 1946 166 0 10 11
0 80 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
969 0 0
2
44771 49
0
13 Logic Switch~
5 2024 163 0 1 11
0 73
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 B3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8402 0 0
2
44771 48
0
13 Logic Switch~
5 2583 1862 0 10 11
0 33 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 B2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3751 0 0
2
44771 47
0
13 Logic Switch~
5 2505 1865 0 10 11
0 40 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4292 0 0
2
44771 46
0
13 Logic Switch~
5 951 1791 0 1 11
0 122
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 A1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6118 0 0
2
44771 1
0
13 Logic Switch~
5 1029 1788 0 10 11
0 115 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 B1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
34 0 0
2
44771 0
0
13 Logic Switch~
5 470 89 0 1 11
0 155
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6357 0 0
2
44771 47
0
13 Logic Switch~
5 392 92 0 10 11
0 162 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 A
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
319 0 0
2
44771 46
0
13 Logic Switch~
5 308 89 0 10 11
0 165 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 Cin
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3976 0 0
2
44771 45
0
13 Logic Switch~
5 234 82 0 1 11
0 4
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 S0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7634 0 0
2
44771 44
0
13 Logic Switch~
5 160 85 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 S1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
523 0 0
2
44771 43
0
13 Logic Switch~
5 82 85 0 1 11
0 6
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 S2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6748 0 0
2
44771 42
0
5 4030~
219 2132 255 0 3 22
0 2 80 90
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U32D
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 32 0
1 U
6901 0 0
2
44771 95
0
9 Inverter~
13 1675 208 0 2 22
0 6 76
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U55F
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 55 0
1 U
842 0 0
2
44771 94
0
9 Inverter~
13 1750 213 0 2 22
0 5 81
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U55E
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 55 0
1 U
3277 0 0
2
44771 93
0
9 Inverter~
13 1824 214 0 2 22
0 4 75
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U55D
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 55 0
1 U
4212 0 0
2
44771 92
0
9 Inverter~
13 1893 212 0 2 22
0 2 74
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U55C
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 55 0
1 U
4720 0 0
2
44771 91
0
9 Inverter~
13 1981 218 0 2 22
0 80 78
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U55B
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 55 0
1 U
5551 0 0
2
44771 90
0
9 Inverter~
13 2064 210 0 2 22
0 73 84
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U55A
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 55 0
1 U
6986 0 0
2
44771 89
0
9 2-In AND~
219 2188 267 0 3 22
0 90 84 89
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U54D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 54 0
1 U
8745 0 0
2
44771 88
0
9 2-In AND~
219 2262 278 0 3 22
0 89 71 62
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U54C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 54 0
1 U
9592 0 0
2
44771 87
0
9 2-In AND~
219 2166 302 0 3 22
0 76 81 71
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U54B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 54 0
1 U
8748 0 0
2
44771 86
0
5 4030~
219 2145 412 0 3 22
0 4 2 88
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U32C
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 32 0
1 U
7168 0 0
2
44771 85
0
5 4030~
219 2193 445 0 3 22
0 88 80 70
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U32B
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 32 0
1 U
631 0 0
2
44771 84
0
9 2-In AND~
219 2204 502 0 3 22
0 76 73 87
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U54A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 54 0
1 U
9466 0 0
2
44771 83
0
9 2-In AND~
219 2273 467 0 3 22
0 70 87 63
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U45D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 45 0
1 U
3266 0 0
2
44771 82
0
5 7415~
219 2205 553 0 4 22
0 76 5 74 66
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U53A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 53 0
1 U
7693 0 0
2
44771 81
0
9 2-In AND~
219 2206 597 0 3 22
0 78 84 65
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U34D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 34 0
1 U
3723 0 0
2
44771 80
0
9 2-In AND~
219 2280 572 0 3 22
0 66 65 64
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U34C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 34 0
1 U
3440 0 0
2
44771 79
0
9 2-In AND~
219 2214 697 0 3 22
0 86 73 61
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U34B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 34 0
1 U
6263 0 0
2
44771 78
0
9 4-In AND~
219 2160 658 0 5 22
0 76 5 4 2 86
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U52B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 52 0
1 U
4900 0 0
2
44771 77
0
9 4-In AND~
219 2167 749 0 5 22
0 5 75 2 80 85
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U52A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 52 0
1 U
8783 0 0
2
44771 76
0
9 2-In AND~
219 2213 787 0 3 22
0 85 84 69
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U45C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 45 0
1 U
3221 0 0
2
44771 75
0
9 4-In AND~
219 2218 844 0 5 22
0 6 5 4 80 83
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U51B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 51 0
1 U
3215 0 0
2
44771 74
0
9 4-In AND~
219 2220 909 0 5 22
0 6 75 78 73 68
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U51A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 51 0
1 U
7903 0 0
2
44771 73
0
9 4-In AND~
219 2220 968 0 5 22
0 174 75 80 84 67
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U50B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 512 2 2 50 0
1 U
7121 0 0
2
44771 72
0
9 4-In AND~
219 2221 1028 0 5 22
0 6 81 78 175 58
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U50A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 512 2 1 50 0
1 U
4484 0 0
2
44771 71
0
8 4-In OR~
219 2350 519 0 5 22
0 62 63 64 61 60
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U49B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 49 0
1 U
5996 0 0
2
44771 70
0
8 4-In OR~
219 2299 844 0 5 22
0 69 83 68 67 59
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U49A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 49 0
1 U
7804 0 0
2
44771 69
0
8 3-In OR~
219 2437 699 0 4 22
0 60 59 58 8
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U44B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 44 0
1 U
5523 0 0
2
44771 68
0
14 Logic Display~
6 2503 624 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3330 0 0
2
44771 67
0
9 4-In AND~
219 2219 1119 0 5 22
0 76 81 2 80 53
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U48B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 48 0
1 U
3465 0 0
2
44771 66
0
9 4-In AND~
219 2223 1193 0 5 22
0 76 81 4 2 82
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U48A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 48 0
1 U
8396 0 0
2
44771 65
0
9 4-In AND~
219 2230 1319 0 5 22
0 76 81 4 80 79
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U47B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 47 0
1 U
3685 0 0
2
44771 64
0
9 4-In AND~
219 2205 1449 0 5 22
0 76 5 74 78 56
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U47A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 47 0
1 U
7849 0 0
2
44771 63
0
9 4-In AND~
219 2229 1549 0 5 22
0 76 5 75 78 77
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U46B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 46 0
1 U
6343 0 0
2
44771 62
0
9 4-In AND~
219 2234 1661 0 5 22
0 76 5 75 74 72
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U46A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 46 0
1 U
7376 0 0
2
44771 61
0
9 2-In AND~
219 2289 1231 0 3 22
0 82 73 52
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U45B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 45 0
1 U
9156 0 0
2
44771 60
0
9 2-In AND~
219 2285 1352 0 3 22
0 79 73 57
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U45A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 45 0
1 U
5776 0 0
2
44771 59
0
9 2-In AND~
219 2313 1591 0 3 22
0 77 73 55
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U42D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 42 0
1 U
7207 0 0
2
44771 58
0
9 2-In AND~
219 2288 1704 0 3 22
0 72 73 54
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U42C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 42 0
1 U
4459 0 0
2
44771 57
0
8 4-In OR~
219 2412 1570 0 5 22
0 57 56 55 54 51
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U43B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 43 0
1 U
3760 0 0
2
44771 56
0
8 3-In OR~
219 2460 1211 0 4 22
0 53 52 51 7
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U44A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 44 0
1 U
754 0 0
2
44771 55
0
14 Logic Display~
6 3104 2867 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9767 0 0
2
44771 41
0
8 3-In OR~
219 3019 2910 0 4 22
0 13 12 11 9
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U21C
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 21 0
1 U
7978 0 0
2
44771 40
0
8 4-In OR~
219 2971 3269 0 5 22
0 17 16 15 14 11
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U43A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 43 0
1 U
3142 0 0
2
44771 39
0
9 2-In AND~
219 2847 3403 0 3 22
0 32 33 14
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U42B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 42 0
1 U
3284 0 0
2
44771 38
0
9 2-In AND~
219 2872 3290 0 3 22
0 37 33 15
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U42A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 42 0
1 U
659 0 0
2
44771 37
0
9 2-In AND~
219 2844 3051 0 3 22
0 39 33 17
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U33D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 33 0
1 U
3800 0 0
2
44771 36
0
9 2-In AND~
219 2848 2930 0 3 22
0 42 33 12
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U33C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 33 0
1 U
6792 0 0
2
44771 35
0
9 4-In AND~
219 2793 3360 0 5 22
0 36 5 35 34 32
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U41B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 41 0
1 U
3701 0 0
2
44771 34
0
9 4-In AND~
219 2788 3248 0 5 22
0 36 5 35 38 37
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U41A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 41 0
1 U
6316 0 0
2
44771 33
0
9 4-In AND~
219 2764 3148 0 5 22
0 36 5 34 38 16
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U40B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 40 0
1 U
8734 0 0
2
44771 32
0
9 4-In AND~
219 2789 3018 0 5 22
0 36 41 4 40 39
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U40A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 40 0
1 U
7988 0 0
2
44771 31
0
9 4-In AND~
219 2782 2892 0 5 22
0 36 41 4 7 42
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U39B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 39 0
1 U
3217 0 0
2
44771 30
0
9 4-In AND~
219 2778 2818 0 5 22
0 36 41 7 40 13
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U39A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 39 0
1 U
3965 0 0
2
44771 29
0
14 Logic Display~
6 3066 2349 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8239 0 0
2
44771 28
0
8 3-In OR~
219 2996 2398 0 4 22
0 20 19 18 10
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U21B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 21 0
1 U
828 0 0
2
44771 27
0
8 4-In OR~
219 2858 2543 0 5 22
0 29 43 28 27 19
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U38B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 38 0
1 U
6187 0 0
2
44771 26
0
8 4-In OR~
219 2909 2218 0 5 22
0 22 23 24 21 20
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U38A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 38 0
1 U
7107 0 0
2
44771 25
0
9 4-In AND~
219 2780 2727 0 5 22
0 6 41 38 176 18
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U37B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 512 2 2 37 0
1 U
6433 0 0
2
44771 24
0
9 4-In AND~
219 2779 2667 0 5 22
0 177 35 40 44 27
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U37A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 512 2 1 37 0
1 U
8559 0 0
2
44771 23
0
9 4-In AND~
219 2779 2608 0 5 22
0 6 35 38 33 28
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U36B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 36 0
1 U
3674 0 0
2
44771 22
0
9 4-In AND~
219 2777 2543 0 5 22
0 6 5 4 40 43
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U36A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 36 0
1 U
5697 0 0
2
44771 21
0
9 2-In AND~
219 2772 2486 0 3 22
0 45 44 29
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U33B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 33 0
1 U
3805 0 0
2
44771 20
0
9 4-In AND~
219 2726 2448 0 5 22
0 5 35 7 40 45
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U35B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 35 0
1 U
5219 0 0
2
44771 19
0
9 4-In AND~
219 2719 2357 0 5 22
0 36 5 4 7 46
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U35A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 35 0
1 U
3795 0 0
2
44771 18
0
9 2-In AND~
219 2773 2396 0 3 22
0 46 33 21
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U34A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 34 0
1 U
3637 0 0
2
44771 17
0
9 2-In AND~
219 2839 2271 0 3 22
0 26 25 24
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U26D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 26 0
1 U
3226 0 0
2
44771 16
0
9 2-In AND~
219 2765 2296 0 3 22
0 38 44 25
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U26C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 26 0
1 U
6966 0 0
2
44771 15
0
5 7415~
219 2764 2252 0 4 22
0 36 5 34 26
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U13C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 13 0
1 U
9796 0 0
2
44771 14
0
9 2-In AND~
219 2832 2166 0 3 22
0 30 47 23
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U33A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 33 0
1 U
5952 0 0
2
44771 13
0
9 2-In AND~
219 2763 2201 0 3 22
0 36 33 47
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U31D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 31 0
1 U
3649 0 0
2
44771 12
0
5 4030~
219 2752 2144 0 3 22
0 48 40 30
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U32A
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 32 0
1 U
3716 0 0
2
44771 11
0
5 4030~
219 2704 2111 0 3 22
0 4 7 48
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U28D
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 28 0
1 U
4797 0 0
2
44771 10
0
9 2-In AND~
219 2725 2001 0 3 22
0 36 41 31
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U31C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 31 0
1 U
4681 0 0
2
44771 9
0
9 2-In AND~
219 2821 1977 0 3 22
0 49 31 22
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U31B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 31 0
1 U
9730 0 0
2
44771 8
0
9 2-In AND~
219 2747 1966 0 3 22
0 50 44 49
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U31A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 31 0
1 U
9874 0 0
2
44771 7
0
9 Inverter~
13 2623 1909 0 2 22
0 33 44
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U30F
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 30 0
1 U
364 0 0
2
44771 6
0
9 Inverter~
13 2540 1917 0 2 22
0 40 38
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U30E
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 30 0
1 U
3656 0 0
2
44771 5
0
9 Inverter~
13 2452 1911 0 2 22
0 7 34
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U30D
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 30 0
1 U
3131 0 0
2
44771 4
0
9 Inverter~
13 2383 1913 0 2 22
0 4 35
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U30C
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 30 0
1 U
6772 0 0
2
44771 3
0
9 Inverter~
13 2309 1912 0 2 22
0 5 41
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U30B
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 30 0
1 U
9557 0 0
2
44771 2
0
9 Inverter~
13 2234 1907 0 2 22
0 6 36
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U30A
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 30 0
1 U
5789 0 0
2
44771 1
0
5 4030~
219 2691 1954 0 3 22
0 7 40 50
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U28C
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 28 0
1 U
7328 0 0
2
44771 0
0
5 4030~
219 1137 1880 0 3 22
0 3 122 132
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U28B
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 28 0
1 U
4799 0 0
2
44771 47
0
9 Inverter~
13 680 1833 0 2 22
0 6 118
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U29F
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 29 0
1 U
9196 0 0
2
44771 46
0
9 Inverter~
13 755 1838 0 2 22
0 5 123
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U29E
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 29 0
1 U
3857 0 0
2
44771 45
0
9 Inverter~
13 829 1839 0 2 22
0 4 117
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U29D
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 29 0
1 U
7125 0 0
2
44771 44
0
9 Inverter~
13 898 1837 0 2 22
0 3 116
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U29C
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 29 0
1 U
3641 0 0
2
44771 43
0
9 Inverter~
13 986 1843 0 2 22
0 122 120
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U29B
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 29 0
1 U
9821 0 0
2
44771 42
0
9 Inverter~
13 1069 1835 0 2 22
0 115 126
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U29A
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 29 0
1 U
3187 0 0
2
44771 41
0
9 2-In AND~
219 1193 1892 0 3 22
0 132 126 131
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U27D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 27 0
1 U
762 0 0
2
44771 40
0
9 2-In AND~
219 1267 1903 0 3 22
0 131 113 104
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U27C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 27 0
1 U
39 0 0
2
44771 39
0
9 2-In AND~
219 1171 1927 0 3 22
0 118 123 113
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U27B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 27 0
1 U
9450 0 0
2
44771 38
0
5 4030~
219 1150 2037 0 3 22
0 4 3 130
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U28A
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 28 0
1 U
3236 0 0
2
44771 37
0
5 4030~
219 1198 2070 0 3 22
0 130 122 112
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U14D
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 14 0
1 U
3321 0 0
2
44771 36
0
9 2-In AND~
219 1209 2127 0 3 22
0 118 115 129
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U27A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 27 0
1 U
8879 0 0
2
44771 35
0
9 2-In AND~
219 1278 2092 0 3 22
0 112 129 105
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U17D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 17 0
1 U
5433 0 0
2
44771 34
0
5 7415~
219 1210 2178 0 4 22
0 118 5 116 108
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U13B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 13 0
1 U
3679 0 0
2
44771 33
0
9 2-In AND~
219 1211 2222 0 3 22
0 120 126 107
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U26B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 26 0
1 U
9342 0 0
2
44771 32
0
9 2-In AND~
219 1285 2197 0 3 22
0 108 107 106
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U26A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 26 0
1 U
3623 0 0
2
44771 31
0
9 2-In AND~
219 1219 2322 0 3 22
0 128 115 103
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U12D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 12 0
1 U
3722 0 0
2
44771 30
0
9 4-In AND~
219 1165 2283 0 5 22
0 118 5 4 3 128
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U25B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 25 0
1 U
8993 0 0
2
44771 29
0
9 4-In AND~
219 1172 2374 0 5 22
0 5 117 3 122 127
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U25A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 25 0
1 U
3723 0 0
2
44771 28
0
9 2-In AND~
219 1218 2412 0 3 22
0 127 126 111
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U17C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 17 0
1 U
6244 0 0
2
44771 27
0
9 4-In AND~
219 1223 2469 0 5 22
0 6 5 4 122 125
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U24B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 24 0
1 U
6421 0 0
2
44771 26
0
9 4-In AND~
219 1225 2534 0 5 22
0 6 117 120 115 110
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U24A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 24 0
1 U
7743 0 0
2
44771 25
0
9 4-In AND~
219 1225 2593 0 5 22
0 178 117 122 126 109
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U23B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 512 2 2 23 0
1 U
9840 0 0
2
44771 24
0
9 4-In AND~
219 1226 2653 0 5 22
0 6 123 120 179 100
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U23A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 512 2 1 23 0
1 U
6910 0 0
2
44771 23
0
8 4-In OR~
219 1355 2144 0 5 22
0 104 105 106 103 102
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U22B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 22 0
1 U
449 0 0
2
44771 22
0
8 4-In OR~
219 1304 2469 0 5 22
0 111 125 110 109 101
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U22A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 22 0
1 U
8761 0 0
2
44771 21
0
8 3-In OR~
219 1442 2324 0 4 22
0 102 101 100 92
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U21A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 21 0
1 U
6748 0 0
2
44771 20
0
14 Logic Display~
6 1512 2275 0 1 2
10 92
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7393 0 0
2
44771 19
0
9 4-In AND~
219 1224 2744 0 5 22
0 118 123 3 122 95
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U20B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 20 0
1 U
7699 0 0
2
44771 18
0
9 4-In AND~
219 1228 2818 0 5 22
0 118 123 4 3 124
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U20A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 20 0
1 U
6638 0 0
2
44771 17
0
9 4-In AND~
219 1235 2944 0 5 22
0 118 123 4 122 121
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U19B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 19 0
1 U
4595 0 0
2
44771 16
0
9 4-In AND~
219 1210 3074 0 5 22
0 118 5 116 120 98
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U19A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 19 0
1 U
9395 0 0
2
44771 15
0
9 4-In AND~
219 1234 3174 0 5 22
0 118 5 117 120 119
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U18B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 18 0
1 U
3303 0 0
2
44771 14
0
9 4-In AND~
219 1239 3286 0 5 22
0 118 5 117 116 114
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U18A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 18 0
1 U
4498 0 0
2
44771 13
0
9 2-In AND~
219 1294 2856 0 3 22
0 124 115 94
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U17B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 17 0
1 U
9728 0 0
2
44771 12
0
9 2-In AND~
219 1290 2977 0 3 22
0 121 115 99
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U17A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 17 0
1 U
3789 0 0
2
44771 11
0
9 2-In AND~
219 1318 3216 0 3 22
0 119 115 97
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U15D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 15 0
1 U
3978 0 0
2
44771 10
0
9 2-In AND~
219 1293 3329 0 3 22
0 114 115 96
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U15C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 15 0
1 U
3494 0 0
2
44771 9
0
8 4-In OR~
219 1417 3195 0 5 22
0 99 98 97 96 93
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U7B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 7 0
1 U
3507 0 0
2
44771 8
0
8 3-In OR~
219 1465 2836 0 4 22
0 95 94 93 2
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U1C
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 1 0
1 U
5151 0 0
2
44771 7
0
8 3-In OR~
219 906 1137 0 4 22
0 135 134 133 3
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U1A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 1 0
1 U
3701 0 0
2
44771 40
0
8 4-In OR~
219 858 1496 0 5 22
0 139 138 137 136 133
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U2A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 2 0
1 U
8585 0 0
2
44771 39
0
9 2-In AND~
219 734 1630 0 3 22
0 154 155 136
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
8809 0 0
2
44771 38
0
9 2-In AND~
219 759 1517 0 3 22
0 159 155 137
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
5993 0 0
2
44771 37
0
9 2-In AND~
219 731 1278 0 3 22
0 161 155 139
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
8654 0 0
2
44771 36
0
9 2-In AND~
219 735 1157 0 3 22
0 164 155 134
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
7223 0 0
2
44771 35
0
9 4-In AND~
219 680 1587 0 5 22
0 158 5 157 156 154
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U4A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 4 0
1 U
3641 0 0
2
44771 34
0
9 4-In AND~
219 675 1475 0 5 22
0 158 5 157 160 159
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U4B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 4 0
1 U
3104 0 0
2
44771 33
0
9 4-In AND~
219 651 1375 0 5 22
0 158 5 156 160 138
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U5A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 5 0
1 U
3296 0 0
2
44771 32
0
9 4-In AND~
219 676 1245 0 5 22
0 158 163 4 162 161
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U5B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 5 0
1 U
8534 0 0
2
44771 31
0
9 4-In AND~
219 669 1119 0 5 22
0 158 163 4 165 164
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U6A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 6 0
1 U
949 0 0
2
44771 30
0
9 4-In AND~
219 665 1045 0 5 22
0 158 163 165 162 135
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U6B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 6 0
1 U
3371 0 0
2
44771 29
0
14 Logic Display~
6 949 550 0 1 2
10 91
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7311 0 0
2
44771 28
0
8 3-In OR~
219 883 625 0 4 22
0 142 141 140 91
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U1B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 1 0
1 U
3409 0 0
2
44771 27
0
8 4-In OR~
219 745 770 0 5 22
0 151 166 150 149 141
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U2B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 2 0
1 U
3526 0 0
2
44771 26
0
8 4-In OR~
219 796 445 0 5 22
0 144 145 146 143 142
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U7A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 7 0
1 U
4129 0 0
2
44771 25
0
9 4-In AND~
219 667 954 0 5 22
0 6 163 160 180 140
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U8A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 512 2 1 8 0
1 U
6278 0 0
2
44771 24
0
9 4-In AND~
219 666 894 0 5 22
0 181 157 162 167 149
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U8B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 512 2 2 8 0
1 U
3482 0 0
2
44771 23
0
9 4-In AND~
219 666 835 0 5 22
0 6 157 160 155 150
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U9A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 9 0
1 U
8323 0 0
2
44771 22
0
9 4-In AND~
219 664 770 0 5 22
0 6 5 4 162 166
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U9B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 9 0
1 U
3984 0 0
2
44771 21
0
9 2-In AND~
219 659 713 0 3 22
0 168 167 151
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U10A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
7622 0 0
2
44771 20
0
9 4-In AND~
219 613 675 0 5 22
0 5 157 165 162 168
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U11A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 11 0
1 U
816 0 0
2
44771 19
0
9 4-In AND~
219 606 584 0 5 22
0 158 5 4 165 169
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U11B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 11 0
1 U
4656 0 0
2
44771 18
0
9 2-In AND~
219 660 623 0 3 22
0 169 155 143
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U12A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
6356 0 0
2
44771 17
0
9 2-In AND~
219 726 498 0 3 22
0 148 147 146
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U12B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 12 0
1 U
7479 0 0
2
44771 16
0
9 2-In AND~
219 652 523 0 3 22
0 160 167 147
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U12C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 12 0
1 U
5690 0 0
2
44771 15
0
5 7415~
219 651 479 0 4 22
0 158 5 156 148
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U13A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 13 0
1 U
5617 0 0
2
44771 14
0
9 2-In AND~
219 719 393 0 3 22
0 152 170 145
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U10B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
3903 0 0
2
44771 13
0
9 2-In AND~
219 650 428 0 3 22
0 158 155 170
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U10C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
4452 0 0
2
44771 12
0
5 4030~
219 639 371 0 3 22
0 171 162 152
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U14A
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 14 0
1 U
6282 0 0
2
44771 11
0
5 4030~
219 591 338 0 3 22
0 4 165 171
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U14B
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 14 0
1 U
7187 0 0
2
44771 10
0
9 2-In AND~
219 612 228 0 3 22
0 158 163 153
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U10D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 10 0
1 U
6866 0 0
2
44771 9
0
9 2-In AND~
219 708 204 0 3 22
0 172 153 144
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U15A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
7670 0 0
2
44771 8
0
9 2-In AND~
219 634 193 0 3 22
0 173 167 172
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U15B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 15 0
1 U
951 0 0
2
44771 7
0
9 Inverter~
13 510 136 0 2 22
0 155 167
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U16A
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 16 0
1 U
9536 0 0
2
44771 6
0
9 Inverter~
13 427 144 0 2 22
0 162 160
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U16B
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 16 0
1 U
5495 0 0
2
44771 5
0
9 Inverter~
13 339 138 0 2 22
0 165 156
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U16C
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 16 0
1 U
8152 0 0
2
44771 4
0
9 Inverter~
13 270 140 0 2 22
0 4 157
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U16D
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 16 0
1 U
6223 0 0
2
44771 3
0
9 Inverter~
13 196 139 0 2 22
0 5 163
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U16E
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 16 0
1 U
5441 0 0
2
44771 2
0
9 Inverter~
13 121 134 0 2 22
0 6 158
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U16F
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 16 0
1 U
3189 0 0
2
44771 1
0
5 4030~
219 578 181 0 3 22
0 165 162 173
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U14C
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 14 0
1 U
8460 0 0
2
44771 0
0
505
0 0 2 0 0 4096 0 0 0 262 13 2
1508 2836
1514 2836
0 0 3 0 0 12288 0 0 0 375 260 4
868 1808
868 1608
968 1608
968 1137
0 0 4 0 0 4096 0 0 0 136 257 2
2343 1980
1783 1980
0 0 5 0 0 4096 0 0 0 137 258 2
2279 1944
1720 1944
0 0 6 0 0 4096 0 0 0 132 259 2
2212 1888
1653 1888
0 0 4 0 0 4096 0 0 0 257 503 4
1784 373
676 373
676 391
229 391
0 0 5 0 0 4096 0 0 0 258 504 2
1720 284
166 284
0 0 6 0 0 4096 0 0 0 259 505 2
1653 218
99 218
0 0 4 0 0 0 0 0 0 382 503 2
789 1914
229 1914
0 0 5 0 0 0 0 0 0 383 504 2
725 1876
166 1876
0 0 6 0 0 0 0 0 0 384 505 2
641 1811
99 1811
0 0 7 0 0 4096 0 0 0 14 135 5
2494 1211
2494 1887
2426 1887
2426 1878
2421 1878
0 0 2 0 0 12304 0 0 0 250 262 6
1862 183
1862 148
1586 148
1586 2758
1514 2758
1514 2836
4 0 7 0 0 0 0 53 0 0 0 3
2493 1211
2523 1211
2523 1144
4 1 8 0 0 8320 0 40 41 0 0 3
2470 699
2503 699
2503 642
4 1 9 0 0 4224 0 55 54 0 0 3
3052 2910
3104 2910
3104 2885
4 1 10 0 0 4224 0 68 67 0 0 3
3029 2398
3066 2398
3066 2367
5 3 11 0 0 8320 0 56 55 0 0 6
3004 3269
3008 3269
3008 2929
3001 2929
3001 2919
3006 2919
3 2 12 0 0 4224 0 60 55 0 0 4
2869 2930
2998 2930
2998 2910
3007 2910
5 1 13 0 0 4224 0 66 55 0 0 4
2799 2818
2998 2818
2998 2901
3006 2901
3 4 14 0 0 8320 0 57 56 0 0 4
2868 3403
2941 3403
2941 3283
2954 3283
3 3 15 0 0 4224 0 58 56 0 0 4
2893 3290
2946 3290
2946 3274
2954 3274
5 2 16 0 0 4224 0 63 56 0 0 4
2785 3148
2941 3148
2941 3265
2954 3265
3 1 17 0 0 8320 0 59 56 0 0 4
2865 3051
2946 3051
2946 3256
2954 3256
5 3 18 0 0 8320 0 71 68 0 0 4
2801 2727
2970 2727
2970 2407
2983 2407
5 2 19 0 0 8320 0 69 68 0 0 4
2891 2543
2975 2543
2975 2398
2984 2398
5 1 20 0 0 8320 0 70 68 0 0 4
2942 2218
2975 2218
2975 2389
2983 2389
3 4 21 0 0 8320 0 78 70 0 0 4
2794 2396
2879 2396
2879 2232
2892 2232
3 1 22 0 0 8320 0 87 70 0 0 4
2842 1977
2879 1977
2879 2205
2892 2205
3 2 23 0 0 8320 0 82 70 0 0 4
2853 2166
2884 2166
2884 2214
2892 2214
3 3 24 0 0 8320 0 79 70 0 0 4
2860 2271
2884 2271
2884 2223
2892 2223
3 2 25 0 0 4224 0 80 79 0 0 4
2786 2296
2807 2296
2807 2280
2815 2280
4 1 26 0 0 4224 0 81 79 0 0 4
2785 2252
2807 2252
2807 2262
2815 2262
5 4 27 0 0 8320 0 72 69 0 0 4
2800 2667
2828 2667
2828 2557
2841 2557
5 3 28 0 0 8320 0 73 69 0 0 4
2800 2608
2833 2608
2833 2548
2841 2548
3 1 29 0 0 8320 0 75 69 0 0 4
2793 2486
2833 2486
2833 2530
2841 2530
3 1 30 0 0 4224 0 84 82 0 0 4
2785 2144
2800 2144
2800 2157
2808 2157
3 2 31 0 0 4224 0 86 87 0 0 4
2746 2001
2789 2001
2789 1986
2797 1986
5 1 32 0 0 8320 0 61 57 0 0 4
2814 3360
2818 3360
2818 3394
2823 3394
2 0 33 0 0 4096 0 57 0 0 133 4
2823 3412
2591 3412
2591 3413
2586 3413
4 0 34 0 0 4096 0 61 0 0 124 2
2769 3374
2456 3374
3 0 35 0 0 4096 0 61 0 0 125 2
2769 3365
2386 3365
2 0 5 0 0 0 0 61 0 0 137 2
2769 3356
2279 3356
1 0 36 0 0 4096 0 61 0 0 122 2
2769 3347
2237 3347
5 1 37 0 0 8320 0 62 58 0 0 4
2809 3248
2840 3248
2840 3281
2848 3281
2 0 33 0 0 4096 0 58 0 0 133 2
2848 3299
2586 3299
4 0 38 0 0 4096 0 62 0 0 123 2
2764 3262
2542 3262
3 0 35 0 0 0 0 62 0 0 125 2
2764 3253
2386 3253
2 0 5 0 0 0 0 62 0 0 137 2
2764 3244
2279 3244
1 0 36 0 0 0 0 62 0 0 122 2
2764 3235
2237 3235
4 0 38 0 0 0 0 63 0 0 123 4
2740 3162
2547 3162
2547 3163
2542 3163
3 0 34 0 0 0 0 63 0 0 124 2
2740 3153
2456 3153
2 0 5 0 0 0 0 63 0 0 137 2
2740 3144
2279 3144
1 0 36 0 0 0 0 63 0 0 122 2
2740 3135
2237 3135
5 1 39 0 0 8320 0 64 59 0 0 4
2810 3018
2814 3018
2814 3042
2820 3042
2 0 33 0 0 0 0 59 0 0 133 2
2820 3060
2586 3060
4 0 40 0 0 4096 0 64 0 0 134 2
2765 3032
2503 3032
3 0 4 0 0 0 0 64 0 0 136 2
2765 3023
2342 3023
2 0 41 0 0 4096 0 64 0 0 126 2
2765 3014
2313 3014
1 0 36 0 0 0 0 64 0 0 122 2
2765 3005
2237 3005
5 1 42 0 0 8320 0 65 60 0 0 4
2803 2892
2816 2892
2816 2921
2824 2921
2 0 33 0 0 0 0 60 0 0 133 2
2824 2939
2586 2939
4 0 7 0 0 0 0 65 0 0 135 2
2758 2906
2417 2906
3 0 4 0 0 0 0 65 0 0 136 2
2758 2897
2342 2897
2 0 41 0 0 0 0 65 0 0 126 2
2758 2888
2313 2888
1 0 36 0 0 0 0 65 0 0 122 2
2758 2879
2237 2879
4 0 40 0 0 0 0 66 0 0 134 2
2754 2832
2503 2832
3 0 7 0 0 0 0 66 0 0 135 2
2754 2823
2417 2823
2 0 41 0 0 0 0 66 0 0 126 2
2754 2814
2313 2814
1 0 36 0 0 0 0 66 0 0 122 2
2754 2805
2237 2805
2 5 43 0 0 4224 0 69 74 0 0 3
2841 2539
2798 2539
2798 2543
0 0 44 0 0 4096 0 0 0 0 119 2
2762 2742
2627 2742
3 0 38 0 0 0 0 71 0 0 123 2
2756 2732
2542 2732
2 0 41 0 0 0 0 71 0 0 126 2
2756 2723
2313 2723
1 0 6 0 0 0 0 71 0 0 138 2
2756 2714
2212 2714
4 0 44 0 0 0 0 72 0 0 119 2
2755 2681
2627 2681
3 0 40 0 0 0 0 72 0 0 134 2
2755 2672
2503 2672
2 0 35 0 0 0 0 72 0 0 125 2
2755 2663
2386 2663
0 0 6 0 0 0 0 0 0 0 138 2
2762 2655
2212 2655
4 0 33 0 0 0 0 73 0 0 133 2
2755 2622
2586 2622
3 0 38 0 0 0 0 73 0 0 123 2
2755 2613
2542 2613
2 0 35 0 0 0 0 73 0 0 125 2
2755 2604
2386 2604
1 0 6 0 0 0 0 73 0 0 138 2
2755 2595
2212 2595
4 0 40 0 0 0 0 74 0 0 134 2
2753 2557
2503 2557
3 0 4 0 0 0 0 74 0 0 136 2
2753 2548
2342 2548
2 0 5 0 0 0 0 74 0 0 137 2
2753 2539
2279 2539
1 0 6 0 0 0 0 74 0 0 138 2
2753 2530
2212 2530
2 0 44 0 0 0 0 75 0 0 119 2
2748 2495
2627 2495
5 1 45 0 0 8320 0 76 75 0 0 3
2747 2448
2748 2448
2748 2477
4 0 40 0 0 0 0 76 0 0 134 2
2702 2462
2503 2462
3 0 7 0 0 0 0 76 0 0 135 2
2702 2453
2417 2453
2 0 35 0 0 0 0 76 0 0 125 2
2702 2444
2386 2444
1 0 5 0 0 0 0 76 0 0 137 2
2702 2435
2279 2435
2 0 33 0 0 0 0 78 0 0 133 2
2749 2405
2586 2405
5 1 46 0 0 8320 0 77 78 0 0 4
2740 2357
2745 2357
2745 2387
2749 2387
4 0 7 0 0 0 0 77 0 0 135 2
2695 2371
2417 2371
3 0 4 0 0 0 0 77 0 0 136 2
2695 2362
2342 2362
2 0 5 0 0 0 0 77 0 0 137 2
2695 2353
2279 2353
1 0 36 0 0 0 0 77 0 0 122 2
2695 2344
2237 2344
2 0 44 0 0 0 0 80 0 0 119 2
2741 2305
2627 2305
1 0 38 0 0 0 0 80 0 0 123 2
2741 2287
2542 2287
3 0 34 0 0 0 0 81 0 0 124 2
2740 2261
2456 2261
2 0 5 0 0 0 0 81 0 0 137 2
2740 2252
2279 2252
1 0 36 0 0 0 0 81 0 0 122 2
2740 2243
2237 2243
2 3 47 0 0 8320 0 82 83 0 0 4
2808 2175
2792 2175
2792 2201
2784 2201
2 0 33 0 0 0 0 83 0 0 133 2
2739 2210
2584 2210
1 0 36 0 0 0 0 83 0 0 122 2
2739 2192
2237 2192
3 1 48 0 0 8320 0 85 84 0 0 4
2737 2111
2728 2111
2728 2135
2736 2135
2 0 40 0 0 0 0 84 0 0 134 2
2736 2153
2503 2153
2 0 7 0 0 0 0 85 0 0 135 4
2688 2120
2422 2120
2422 2123
2417 2123
1 0 4 0 0 0 0 85 0 0 136 4
2688 2102
2358 2102
2358 2104
2343 2104
3 1 49 0 0 8320 0 88 87 0 0 3
2768 1966
2768 1968
2797 1968
2 0 44 0 0 0 0 88 0 0 119 4
2723 1975
2642 1975
2642 1987
2627 1987
3 1 50 0 0 8320 0 95 88 0 0 3
2724 1954
2723 1954
2723 1957
0 2 41 0 0 0 0 0 86 126 0 4
2313 2054
2328 2054
2328 2010
2701 2010
1 0 36 0 0 0 0 86 0 0 122 4
2701 1992
2252 1992
2252 2036
2237 2036
2 0 40 0 0 0 0 95 0 0 134 2
2675 1963
2503 1963
1 0 7 0 0 0 0 95 0 0 135 2
2675 1945
2417 1945
0 2 44 0 0 8320 0 0 89 0 0 4
2628 5245
2627 5245
2627 1927
2626 1927
2 0 38 0 0 0 0 90 0 0 123 3
2543 1935
2548 1935
2548 1930
2 0 34 0 0 0 0 91 0 0 124 4
2455 1929
2455 1926
2455 1926
2455 1939
0 2 36 0 0 8320 0 0 94 0 0 3
2249 5235
2237 5235
2237 1925
0 1 38 0 0 4224 0 0 0 0 0 4
2542 5243
2542 1935
2548 1935
2548 1927
1 0 34 0 0 12416 0 0 0 121 0 4
2455 1926
2455 1939
2456 1939
2456 5241
2 0 35 0 0 4224 0 92 0 0 0 3
2386 1931
2386 5241
2382 5241
2 0 41 0 0 8320 0 93 0 0 0 3
2312 1930
2313 1930
2313 5236
1 0 33 0 0 0 0 89 0 0 133 3
2626 1891
2626 1879
2583 1879
1 0 40 0 0 0 0 90 0 0 134 5
2543 1899
2543 1882
2508 1882
2508 1889
2503 1889
1 0 7 0 0 0 0 91 0 0 135 3
2455 1893
2455 1882
2421 1882
1 0 4 0 0 0 0 92 0 0 136 3
2386 1895
2386 1882
2343 1882
1 0 5 0 0 0 0 93 0 0 137 3
2312 1894
2312 1882
2278 1882
1 0 6 0 0 0 0 94 0 0 138 5
2237 1889
2237 1883
2212 1883
2212 1888
2207 1888
1 0 33 0 0 20608 0 3 0 0 0 6
2583 1874
2583 1924
2584 1924
2584 2210
2586 2210
2586 5217
0 1 40 0 0 8320 0 0 4 0 0 5
2502 5213
2503 5213
2503 1885
2505 1885
2505 1877
0 0 7 0 0 12416 0 0 0 0 0 5
2421 1874
2421 1889
2417 1889
2417 5211
2418 5211
0 0 4 0 0 16512 0 0 0 0 0 5
2347 1867
2343 1867
2343 2104
2342 2104
2342 5211
0 0 5 0 0 16512 0 0 0 0 0 5
2273 1870
2278 1870
2278 1921
2279 1921
2279 5209
0 0 6 0 0 20608 0 0 0 0 0 6
2195 1870
2195 1885
2207 1885
2207 1888
2212 1888
2212 5206
5 3 51 0 0 8320 0 52 53 0 0 6
2445 1570
2449 1570
2449 1230
2442 1230
2442 1220
2447 1220
3 2 52 0 0 4224 0 48 53 0 0 4
2310 1231
2439 1231
2439 1211
2448 1211
5 1 53 0 0 4224 0 42 53 0 0 4
2240 1119
2439 1119
2439 1202
2447 1202
3 4 54 0 0 8320 0 51 52 0 0 4
2309 1704
2382 1704
2382 1584
2395 1584
3 3 55 0 0 4224 0 50 52 0 0 4
2334 1591
2387 1591
2387 1575
2395 1575
5 2 56 0 0 4224 0 45 52 0 0 4
2226 1449
2382 1449
2382 1566
2395 1566
3 1 57 0 0 8320 0 49 52 0 0 4
2306 1352
2387 1352
2387 1557
2395 1557
5 3 58 0 0 8320 0 37 40 0 0 4
2242 1028
2411 1028
2411 708
2424 708
5 2 59 0 0 8320 0 39 40 0 0 4
2332 844
2416 844
2416 699
2425 699
5 1 60 0 0 8320 0 38 40 0 0 4
2383 519
2416 519
2416 690
2424 690
3 4 61 0 0 8320 0 30 38 0 0 4
2235 697
2320 697
2320 533
2333 533
3 1 62 0 0 8320 0 21 38 0 0 4
2283 278
2320 278
2320 506
2333 506
3 2 63 0 0 8320 0 26 38 0 0 4
2294 467
2325 467
2325 515
2333 515
3 3 64 0 0 8320 0 29 38 0 0 4
2301 572
2325 572
2325 524
2333 524
3 2 65 0 0 4224 0 28 29 0 0 4
2227 597
2248 597
2248 581
2256 581
4 1 66 0 0 4224 0 27 29 0 0 4
2226 553
2248 553
2248 563
2256 563
5 4 67 0 0 8320 0 36 39 0 0 4
2241 968
2269 968
2269 858
2282 858
5 3 68 0 0 8320 0 35 39 0 0 4
2241 909
2274 909
2274 849
2282 849
3 1 69 0 0 8320 0 33 39 0 0 4
2234 787
2274 787
2274 831
2282 831
3 1 70 0 0 4224 0 24 26 0 0 4
2226 445
2241 445
2241 458
2249 458
3 2 71 0 0 4224 0 22 21 0 0 4
2187 302
2230 302
2230 287
2238 287
5 1 72 0 0 8320 0 47 51 0 0 4
2255 1661
2259 1661
2259 1695
2264 1695
2 0 73 0 0 4096 0 51 0 0 254 4
2264 1713
2032 1713
2032 1714
2027 1714
4 0 74 0 0 4096 0 47 0 0 245 2
2210 1675
1897 1675
3 0 75 0 0 4096 0 47 0 0 246 2
2210 1666
1827 1666
2 0 5 0 0 0 0 47 0 0 258 2
2210 1657
1720 1657
1 0 76 0 0 4096 0 47 0 0 243 2
2210 1648
1678 1648
5 1 77 0 0 8320 0 46 50 0 0 4
2250 1549
2281 1549
2281 1582
2289 1582
2 0 73 0 0 4096 0 50 0 0 254 2
2289 1600
2027 1600
4 0 78 0 0 4096 0 46 0 0 244 2
2205 1563
1983 1563
3 0 75 0 0 0 0 46 0 0 246 2
2205 1554
1827 1554
2 0 5 0 0 0 0 46 0 0 258 2
2205 1545
1720 1545
1 0 76 0 0 0 0 46 0 0 243 2
2205 1536
1678 1536
4 0 78 0 0 0 0 45 0 0 244 4
2181 1463
1988 1463
1988 1464
1983 1464
3 0 74 0 0 0 0 45 0 0 245 2
2181 1454
1897 1454
2 0 5 0 0 0 0 45 0 0 258 2
2181 1445
1720 1445
1 0 76 0 0 0 0 45 0 0 243 2
2181 1436
1678 1436
5 1 79 0 0 8320 0 44 49 0 0 4
2251 1319
2255 1319
2255 1343
2261 1343
2 0 73 0 0 0 0 49 0 0 254 2
2261 1361
2027 1361
4 0 80 0 0 4096 0 44 0 0 255 2
2206 1333
1944 1333
3 0 4 0 0 0 0 44 0 0 257 2
2206 1324
1783 1324
2 0 81 0 0 4096 0 44 0 0 247 2
2206 1315
1754 1315
1 0 76 0 0 0 0 44 0 0 243 2
2206 1306
1678 1306
5 1 82 0 0 8320 0 43 48 0 0 4
2244 1193
2257 1193
2257 1222
2265 1222
2 0 73 0 0 0 0 48 0 0 254 2
2265 1240
2027 1240
4 0 2 0 0 0 0 43 0 0 256 2
2199 1207
1858 1207
3 0 4 0 0 0 0 43 0 0 257 2
2199 1198
1783 1198
2 0 81 0 0 0 0 43 0 0 247 2
2199 1189
1754 1189
1 0 76 0 0 0 0 43 0 0 243 2
2199 1180
1678 1180
4 0 80 0 0 0 0 42 0 0 255 2
2195 1133
1944 1133
3 0 2 0 0 0 0 42 0 0 256 2
2195 1124
1858 1124
2 0 81 0 0 0 0 42 0 0 247 2
2195 1115
1754 1115
1 0 76 0 0 0 0 42 0 0 243 2
2195 1106
1678 1106
2 5 83 0 0 4224 0 39 34 0 0 3
2282 840
2239 840
2239 844
0 0 84 0 0 4096 0 0 0 0 240 2
2203 1043
2068 1043
3 0 78 0 0 0 0 37 0 0 244 2
2197 1033
1983 1033
2 0 81 0 0 0 0 37 0 0 247 2
2197 1024
1754 1024
1 0 6 0 0 0 0 37 0 0 259 2
2197 1015
1653 1015
4 0 84 0 0 0 0 36 0 0 240 2
2196 982
2068 982
3 0 80 0 0 0 0 36 0 0 255 2
2196 973
1944 973
2 0 75 0 0 0 0 36 0 0 246 2
2196 964
1827 964
0 0 6 0 0 0 0 0 0 0 259 2
2203 956
1653 956
4 0 73 0 0 0 0 35 0 0 254 2
2196 923
2027 923
3 0 78 0 0 0 0 35 0 0 244 2
2196 914
1983 914
2 0 75 0 0 0 0 35 0 0 246 2
2196 905
1827 905
1 0 6 0 0 0 0 35 0 0 259 2
2196 896
1653 896
4 0 80 0 0 0 0 34 0 0 255 2
2194 858
1944 858
3 0 4 0 0 0 0 34 0 0 257 2
2194 849
1783 849
2 0 5 0 0 0 0 34 0 0 258 2
2194 840
1720 840
1 0 6 0 0 0 0 34 0 0 259 2
2194 831
1653 831
2 0 84 0 0 0 0 33 0 0 240 2
2189 796
2068 796
5 1 85 0 0 8320 0 32 33 0 0 3
2188 749
2189 749
2189 778
4 0 80 0 0 0 0 32 0 0 255 2
2143 763
1944 763
3 0 2 0 0 0 0 32 0 0 256 2
2143 754
1858 754
2 0 75 0 0 0 0 32 0 0 246 2
2143 745
1827 745
1 0 5 0 0 0 0 32 0 0 258 2
2143 736
1720 736
2 0 73 0 0 0 0 30 0 0 254 2
2190 706
2027 706
5 1 86 0 0 8320 0 31 30 0 0 4
2181 658
2186 658
2186 688
2190 688
4 0 2 0 0 0 0 31 0 0 256 2
2136 672
1858 672
3 0 4 0 0 0 0 31 0 0 257 2
2136 663
1783 663
2 0 5 0 0 0 0 31 0 0 258 2
2136 654
1720 654
1 0 76 0 0 0 0 31 0 0 243 2
2136 645
1678 645
2 0 84 0 0 0 0 28 0 0 240 2
2182 606
2068 606
1 0 78 0 0 0 0 28 0 0 244 2
2182 588
1983 588
3 0 74 0 0 0 0 27 0 0 245 2
2181 562
1897 562
2 0 5 0 0 0 0 27 0 0 258 2
2181 553
1720 553
1 0 76 0 0 0 0 27 0 0 243 2
2181 544
1678 544
2 3 87 0 0 8320 0 26 25 0 0 4
2249 476
2233 476
2233 502
2225 502
2 0 73 0 0 0 0 25 0 0 254 2
2180 511
2025 511
1 0 76 0 0 0 0 25 0 0 243 2
2180 493
1678 493
3 1 88 0 0 8320 0 23 24 0 0 4
2178 412
2169 412
2169 436
2177 436
2 0 80 0 0 0 0 24 0 0 255 2
2177 454
1944 454
2 0 2 0 0 0 0 23 0 0 256 4
2129 421
1863 421
1863 424
1858 424
1 0 4 0 0 0 0 23 0 0 257 4
2129 403
1799 403
1799 405
1784 405
3 1 89 0 0 8320 0 20 21 0 0 3
2209 267
2209 269
2238 269
2 0 84 0 0 0 0 20 0 0 240 4
2164 276
2083 276
2083 288
2068 288
3 1 90 0 0 8320 0 13 20 0 0 3
2165 255
2164 255
2164 258
0 2 81 0 0 0 0 0 22 247 0 4
1754 355
1769 355
1769 311
2142 311
1 0 76 0 0 0 0 22 0 0 243 4
2142 293
1693 293
1693 337
1678 337
2 0 80 0 0 0 0 13 0 0 255 2
2116 264
1944 264
1 0 2 0 0 0 0 13 0 0 256 2
2116 246
1858 246
0 2 84 0 0 8320 0 0 19 0 0 4
2069 3546
2068 3546
2068 228
2067 228
2 0 78 0 0 0 0 18 0 0 244 3
1984 236
1989 236
1989 231
2 0 74 0 0 0 0 17 0 0 245 4
1896 230
1896 227
1896 227
1896 240
0 2 76 0 0 8320 0 0 14 0 0 3
1690 3536
1678 3536
1678 226
0 1 78 0 0 4224 0 0 0 0 0 4
1983 3544
1983 236
1989 236
1989 228
1 0 74 0 0 12416 0 0 0 242 0 4
1896 227
1896 240
1897 240
1897 3542
2 0 75 0 0 4224 0 16 0 0 0 3
1827 232
1827 3542
1823 3542
2 0 81 0 0 8320 0 15 0 0 0 3
1753 231
1754 231
1754 3537
1 0 73 0 0 0 0 19 0 0 254 3
2067 192
2067 180
2024 180
1 0 80 0 0 0 0 18 0 0 255 5
1984 200
1984 183
1949 183
1949 190
1944 190
1 0 2 0 0 0 0 17 0 0 256 3
1896 194
1896 183
1862 183
1 0 4 0 0 0 0 16 0 0 257 3
1827 196
1827 183
1784 183
1 0 5 0 0 0 0 15 0 0 258 3
1753 195
1753 183
1719 183
1 0 6 0 0 0 0 14 0 0 259 5
1678 190
1678 184
1653 184
1653 189
1648 189
1 0 73 0 0 20608 0 2 0 0 0 6
2024 175
2024 225
2025 225
2025 511
2027 511
2027 3518
0 1 80 0 0 8320 0 0 1 0 0 5
1943 3514
1944 3514
1944 186
1946 186
1946 178
0 0 2 0 0 12416 0 0 0 13 0 5
1862 175
1862 190
1858 190
1858 3512
1859 3512
0 0 4 0 0 0 0 0 0 0 0 5
1788 168
1784 168
1784 405
1783 405
1783 3512
0 0 5 0 0 0 0 0 0 0 0 5
1714 171
1719 171
1719 222
1720 222
1720 3510
0 0 6 0 0 0 0 0 0 0 0 6
1636 171
1636 186
1648 186
1648 189
1653 189
1653 3507
4 0 3 0 0 0 0 137 0 0 0 3
939 1137
969 1137
969 1070
4 1 91 0 0 8320 0 150 149 0 0 3
916 625
949 625
949 568
4 0 2 0 0 0 0 136 0 0 0 3
1498 2836
1550 2836
1550 2811
4 1 92 0 0 4224 0 123 124 0 0 3
1475 2324
1512 2324
1512 2293
5 3 93 0 0 8320 0 135 136 0 0 6
1450 3195
1454 3195
1454 2855
1447 2855
1447 2845
1452 2845
3 2 94 0 0 4224 0 131 136 0 0 4
1315 2856
1444 2856
1444 2836
1453 2836
5 1 95 0 0 4224 0 125 136 0 0 4
1245 2744
1444 2744
1444 2827
1452 2827
3 4 96 0 0 8320 0 134 135 0 0 4
1314 3329
1387 3329
1387 3209
1400 3209
3 3 97 0 0 4224 0 133 135 0 0 4
1339 3216
1392 3216
1392 3200
1400 3200
5 2 98 0 0 4224 0 128 135 0 0 4
1231 3074
1387 3074
1387 3191
1400 3191
3 1 99 0 0 8320 0 132 135 0 0 4
1311 2977
1392 2977
1392 3182
1400 3182
5 3 100 0 0 8320 0 120 123 0 0 4
1247 2653
1416 2653
1416 2333
1429 2333
5 2 101 0 0 8320 0 122 123 0 0 4
1337 2469
1421 2469
1421 2324
1430 2324
5 1 102 0 0 8320 0 121 123 0 0 4
1388 2144
1421 2144
1421 2315
1429 2315
3 4 103 0 0 8320 0 113 121 0 0 4
1240 2322
1325 2322
1325 2158
1338 2158
3 1 104 0 0 8320 0 104 121 0 0 4
1288 1903
1325 1903
1325 2131
1338 2131
3 2 105 0 0 8320 0 109 121 0 0 4
1299 2092
1330 2092
1330 2140
1338 2140
3 3 106 0 0 8320 0 112 121 0 0 4
1306 2197
1330 2197
1330 2149
1338 2149
3 2 107 0 0 4224 0 111 112 0 0 4
1232 2222
1253 2222
1253 2206
1261 2206
4 1 108 0 0 4224 0 110 112 0 0 4
1231 2178
1253 2178
1253 2188
1261 2188
5 4 109 0 0 8320 0 119 122 0 0 4
1246 2593
1274 2593
1274 2483
1287 2483
5 3 110 0 0 8320 0 118 122 0 0 4
1246 2534
1279 2534
1279 2474
1287 2474
3 1 111 0 0 8320 0 116 122 0 0 4
1239 2412
1279 2412
1279 2456
1287 2456
3 1 112 0 0 4224 0 107 109 0 0 4
1231 2070
1246 2070
1246 2083
1254 2083
3 2 113 0 0 4224 0 105 104 0 0 4
1192 1927
1235 1927
1235 1912
1243 1912
5 1 114 0 0 8320 0 130 134 0 0 4
1260 3286
1264 3286
1264 3320
1269 3320
2 0 115 0 0 4096 0 134 0 0 379 4
1269 3338
1037 3338
1037 3339
1032 3339
4 0 116 0 0 4096 0 130 0 0 370 2
1215 3300
902 3300
3 0 117 0 0 4096 0 130 0 0 371 2
1215 3291
832 3291
2 0 5 0 0 0 0 130 0 0 383 2
1215 3282
725 3282
1 0 118 0 0 4096 0 130 0 0 368 2
1215 3273
683 3273
5 1 119 0 0 8320 0 129 133 0 0 4
1255 3174
1286 3174
1286 3207
1294 3207
2 0 115 0 0 4096 0 133 0 0 379 2
1294 3225
1032 3225
4 0 120 0 0 4096 0 129 0 0 369 2
1210 3188
988 3188
3 0 117 0 0 0 0 129 0 0 371 2
1210 3179
832 3179
2 0 5 0 0 0 0 129 0 0 383 2
1210 3170
725 3170
1 0 118 0 0 0 0 129 0 0 368 2
1210 3161
683 3161
4 0 120 0 0 0 0 128 0 0 369 4
1186 3088
993 3088
993 3089
988 3089
3 0 116 0 0 0 0 128 0 0 370 2
1186 3079
902 3079
2 0 5 0 0 0 0 128 0 0 383 2
1186 3070
725 3070
1 0 118 0 0 0 0 128 0 0 368 2
1186 3061
683 3061
5 1 121 0 0 8320 0 127 132 0 0 4
1256 2944
1260 2944
1260 2968
1266 2968
2 0 115 0 0 0 0 132 0 0 379 2
1266 2986
1032 2986
4 0 122 0 0 4096 0 127 0 0 380 2
1211 2958
949 2958
3 0 4 0 0 0 0 127 0 0 382 2
1211 2949
788 2949
2 0 123 0 0 4096 0 127 0 0 372 2
1211 2940
759 2940
1 0 118 0 0 0 0 127 0 0 368 2
1211 2931
683 2931
5 1 124 0 0 8320 0 126 131 0 0 4
1249 2818
1262 2818
1262 2847
1270 2847
2 0 115 0 0 0 0 131 0 0 379 2
1270 2865
1032 2865
4 0 3 0 0 0 0 126 0 0 381 2
1204 2832
863 2832
3 0 4 0 0 0 0 126 0 0 382 2
1204 2823
788 2823
2 0 123 0 0 0 0 126 0 0 372 2
1204 2814
759 2814
1 0 118 0 0 0 0 126 0 0 368 2
1204 2805
683 2805
4 0 122 0 0 0 0 125 0 0 380 2
1200 2758
949 2758
3 0 3 0 0 0 0 125 0 0 381 2
1200 2749
863 2749
2 0 123 0 0 0 0 125 0 0 372 2
1200 2740
759 2740
1 0 118 0 0 0 0 125 0 0 368 2
1200 2731
683 2731
2 5 125 0 0 4224 0 122 117 0 0 3
1287 2465
1244 2465
1244 2469
0 0 126 0 0 4096 0 0 0 0 365 2
1208 2668
1073 2668
3 0 120 0 0 0 0 120 0 0 369 2
1202 2658
988 2658
2 0 123 0 0 0 0 120 0 0 372 2
1202 2649
759 2649
1 0 6 0 0 0 0 120 0 0 384 2
1202 2640
658 2640
4 0 126 0 0 0 0 119 0 0 365 2
1201 2607
1073 2607
3 0 122 0 0 0 0 119 0 0 380 2
1201 2598
949 2598
2 0 117 0 0 0 0 119 0 0 371 2
1201 2589
832 2589
0 0 6 0 0 0 0 0 0 0 384 2
1208 2581
658 2581
4 0 115 0 0 0 0 118 0 0 379 2
1201 2548
1032 2548
3 0 120 0 0 0 0 118 0 0 369 2
1201 2539
988 2539
2 0 117 0 0 0 0 118 0 0 371 2
1201 2530
832 2530
1 0 6 0 0 0 0 118 0 0 384 2
1201 2521
658 2521
4 0 122 0 0 0 0 117 0 0 380 2
1199 2483
949 2483
3 0 4 0 0 0 0 117 0 0 382 2
1199 2474
788 2474
2 0 5 0 0 0 0 117 0 0 383 2
1199 2465
725 2465
1 0 6 0 0 0 0 117 0 0 384 2
1199 2456
658 2456
2 0 126 0 0 0 0 116 0 0 365 2
1194 2421
1073 2421
5 1 127 0 0 8320 0 115 116 0 0 3
1193 2374
1194 2374
1194 2403
4 0 122 0 0 0 0 115 0 0 380 2
1148 2388
949 2388
3 0 3 0 0 0 0 115 0 0 381 2
1148 2379
863 2379
2 0 117 0 0 0 0 115 0 0 371 2
1148 2370
832 2370
1 0 5 0 0 0 0 115 0 0 383 2
1148 2361
725 2361
2 0 115 0 0 0 0 113 0 0 379 2
1195 2331
1032 2331
5 1 128 0 0 8320 0 114 113 0 0 4
1186 2283
1191 2283
1191 2313
1195 2313
4 0 3 0 0 0 0 114 0 0 381 2
1141 2297
863 2297
3 0 4 0 0 0 0 114 0 0 382 2
1141 2288
788 2288
2 0 5 0 0 0 0 114 0 0 383 2
1141 2279
725 2279
1 0 118 0 0 0 0 114 0 0 368 2
1141 2270
683 2270
2 0 126 0 0 0 0 111 0 0 365 2
1187 2231
1073 2231
1 0 120 0 0 0 0 111 0 0 369 2
1187 2213
988 2213
3 0 116 0 0 0 0 110 0 0 370 2
1186 2187
902 2187
2 0 5 0 0 0 0 110 0 0 383 2
1186 2178
725 2178
1 0 118 0 0 0 0 110 0 0 368 2
1186 2169
683 2169
2 3 129 0 0 8320 0 109 108 0 0 4
1254 2101
1238 2101
1238 2127
1230 2127
2 0 115 0 0 0 0 108 0 0 379 2
1185 2136
1030 2136
1 0 118 0 0 0 0 108 0 0 368 2
1185 2118
683 2118
3 1 130 0 0 8320 0 106 107 0 0 4
1183 2037
1174 2037
1174 2061
1182 2061
2 0 122 0 0 0 0 107 0 0 380 2
1182 2079
949 2079
2 0 3 0 0 0 0 106 0 0 381 4
1134 2046
868 2046
868 2049
863 2049
1 0 4 0 0 0 0 106 0 0 382 4
1134 2028
804 2028
804 2030
789 2030
3 1 131 0 0 8320 0 103 104 0 0 3
1214 1892
1214 1894
1243 1894
2 0 126 0 0 0 0 103 0 0 365 4
1169 1901
1088 1901
1088 1913
1073 1913
3 1 132 0 0 8320 0 96 103 0 0 3
1170 1880
1169 1880
1169 1883
0 2 123 0 0 0 0 0 105 372 0 4
759 1980
774 1980
774 1936
1147 1936
1 0 118 0 0 0 0 105 0 0 368 4
1147 1918
698 1918
698 1962
683 1962
2 0 122 0 0 0 0 96 0 0 380 2
1121 1889
949 1889
1 0 3 0 0 0 0 96 0 0 381 2
1121 1871
863 1871
0 2 126 0 0 8320 0 0 102 0 0 4
1074 5171
1073 5171
1073 1853
1072 1853
2 0 120 0 0 0 0 101 0 0 369 3
989 1861
994 1861
994 1856
2 0 116 0 0 0 0 100 0 0 370 4
901 1855
901 1852
901 1852
901 1865
0 2 118 0 0 8320 0 0 97 0 0 3
695 5161
683 5161
683 1851
0 1 120 0 0 4224 0 0 0 0 0 4
988 5169
988 1861
994 1861
994 1853
1 0 116 0 0 12416 0 0 0 367 0 4
901 1852
901 1865
902 1865
902 5167
2 0 117 0 0 4224 0 99 0 0 0 3
832 1857
832 5167
828 5167
2 0 123 0 0 8320 0 98 0 0 0 3
758 1856
759 1856
759 5162
1 0 115 0 0 0 0 102 0 0 379 3
1072 1817
1072 1805
1029 1805
1 0 122 0 0 0 0 101 0 0 380 5
989 1825
989 1808
954 1808
954 1815
949 1815
1 0 3 0 0 0 0 100 0 0 381 3
901 1819
901 1808
867 1808
1 0 4 0 0 0 0 99 0 0 382 3
832 1821
832 1808
789 1808
1 0 5 0 0 0 0 98 0 0 383 3
758 1820
758 1808
724 1808
1 0 6 0 0 0 0 97 0 0 384 5
683 1815
683 1809
658 1809
658 1814
653 1814
1 0 115 0 0 20608 0 6 0 0 0 6
1029 1800
1029 1850
1030 1850
1030 2136
1032 2136
1032 5143
0 1 122 0 0 8320 0 0 5 0 0 5
948 5139
949 5139
949 1811
951 1811
951 1803
0 0 3 0 0 12416 0 0 0 0 0 5
867 1800
867 1815
863 1815
863 5137
864 5137
0 0 4 0 0 0 0 0 0 0 0 5
793 1793
789 1793
789 2030
788 2030
788 5137
0 0 5 0 0 0 0 0 0 0 0 5
719 1796
724 1796
724 1847
725 1847
725 5135
0 0 6 0 0 0 0 0 0 0 0 6
641 1796
641 1811
653 1811
653 1814
658 1814
658 5132
5 3 133 0 0 8320 0 138 137 0 0 6
891 1496
895 1496
895 1156
888 1156
888 1146
893 1146
3 2 134 0 0 4224 0 142 137 0 0 4
756 1157
885 1157
885 1137
894 1137
5 1 135 0 0 4224 0 148 137 0 0 4
686 1045
885 1045
885 1128
893 1128
3 4 136 0 0 8320 0 139 138 0 0 4
755 1630
828 1630
828 1510
841 1510
3 3 137 0 0 4224 0 140 138 0 0 4
780 1517
833 1517
833 1501
841 1501
5 2 138 0 0 4224 0 145 138 0 0 4
672 1375
828 1375
828 1492
841 1492
3 1 139 0 0 8320 0 141 138 0 0 4
752 1278
833 1278
833 1483
841 1483
5 3 140 0 0 8320 0 153 150 0 0 4
688 954
857 954
857 634
870 634
5 2 141 0 0 8320 0 151 150 0 0 4
778 770
862 770
862 625
871 625
5 1 142 0 0 8320 0 152 150 0 0 4
829 445
862 445
862 616
870 616
3 4 143 0 0 8320 0 160 152 0 0 4
681 623
766 623
766 459
779 459
3 1 144 0 0 8320 0 169 152 0 0 4
729 204
766 204
766 432
779 432
3 2 145 0 0 8320 0 164 152 0 0 4
740 393
771 393
771 441
779 441
3 3 146 0 0 8320 0 161 152 0 0 4
747 498
771 498
771 450
779 450
3 2 147 0 0 4224 0 162 161 0 0 4
673 523
694 523
694 507
702 507
4 1 148 0 0 4224 0 163 161 0 0 4
672 479
694 479
694 489
702 489
5 4 149 0 0 8320 0 154 151 0 0 4
687 894
715 894
715 784
728 784
5 3 150 0 0 8320 0 155 151 0 0 4
687 835
720 835
720 775
728 775
3 1 151 0 0 8320 0 157 151 0 0 4
680 713
720 713
720 757
728 757
3 1 152 0 0 4224 0 166 164 0 0 4
672 371
687 371
687 384
695 384
3 2 153 0 0 4224 0 168 169 0 0 4
633 228
676 228
676 213
684 213
5 1 154 0 0 8320 0 143 139 0 0 4
701 1587
705 1587
705 1621
710 1621
2 0 155 0 0 4096 0 139 0 0 500 4
710 1639
478 1639
478 1640
473 1640
4 0 156 0 0 4096 0 143 0 0 491 2
656 1601
343 1601
3 0 157 0 0 4096 0 143 0 0 492 2
656 1592
273 1592
2 0 5 0 0 0 0 143 0 0 504 2
656 1583
166 1583
1 0 158 0 0 4096 0 143 0 0 489 2
656 1574
124 1574
5 1 159 0 0 8320 0 144 140 0 0 4
696 1475
727 1475
727 1508
735 1508
2 0 155 0 0 4096 0 140 0 0 500 2
735 1526
473 1526
4 0 160 0 0 4096 0 144 0 0 490 2
651 1489
429 1489
3 0 157 0 0 0 0 144 0 0 492 2
651 1480
273 1480
2 0 5 0 0 0 0 144 0 0 504 2
651 1471
166 1471
1 0 158 0 0 0 0 144 0 0 489 2
651 1462
124 1462
4 0 160 0 0 0 0 145 0 0 490 4
627 1389
434 1389
434 1390
429 1390
3 0 156 0 0 0 0 145 0 0 491 2
627 1380
343 1380
2 0 5 0 0 0 0 145 0 0 504 2
627 1371
166 1371
1 0 158 0 0 0 0 145 0 0 489 2
627 1362
124 1362
5 1 161 0 0 8320 0 146 141 0 0 4
697 1245
701 1245
701 1269
707 1269
2 0 155 0 0 0 0 141 0 0 500 2
707 1287
473 1287
4 0 162 0 0 4096 0 146 0 0 501 2
652 1259
390 1259
3 0 4 0 0 0 0 146 0 0 503 2
652 1250
229 1250
2 0 163 0 0 4096 0 146 0 0 493 2
652 1241
200 1241
1 0 158 0 0 0 0 146 0 0 489 2
652 1232
124 1232
5 1 164 0 0 8320 0 147 142 0 0 4
690 1119
703 1119
703 1148
711 1148
2 0 155 0 0 0 0 142 0 0 500 2
711 1166
473 1166
4 0 165 0 0 4096 0 147 0 0 502 2
645 1133
304 1133
3 0 4 0 0 0 0 147 0 0 503 2
645 1124
229 1124
2 0 163 0 0 0 0 147 0 0 493 2
645 1115
200 1115
1 0 158 0 0 0 0 147 0 0 489 2
645 1106
124 1106
4 0 162 0 0 0 0 148 0 0 501 2
641 1059
390 1059
3 0 165 0 0 0 0 148 0 0 502 2
641 1050
304 1050
2 0 163 0 0 0 0 148 0 0 493 2
641 1041
200 1041
1 0 158 0 0 0 0 148 0 0 489 2
641 1032
124 1032
2 5 166 0 0 4224 0 151 156 0 0 3
728 766
685 766
685 770
0 0 167 0 0 4096 0 0 0 0 486 2
649 969
514 969
3 0 160 0 0 0 0 153 0 0 490 2
643 959
429 959
2 0 163 0 0 0 0 153 0 0 493 2
643 950
200 950
1 0 6 0 0 0 0 153 0 0 505 2
643 941
99 941
4 0 167 0 0 0 0 154 0 0 486 2
642 908
514 908
3 0 162 0 0 0 0 154 0 0 501 2
642 899
390 899
2 0 157 0 0 0 0 154 0 0 492 2
642 890
273 890
0 0 6 0 0 0 0 0 0 0 505 2
649 882
99 882
4 0 155 0 0 0 0 155 0 0 500 2
642 849
473 849
3 0 160 0 0 0 0 155 0 0 490 2
642 840
429 840
2 0 157 0 0 0 0 155 0 0 492 2
642 831
273 831
1 0 6 0 0 0 0 155 0 0 505 2
642 822
99 822
4 0 162 0 0 0 0 156 0 0 501 2
640 784
390 784
3 0 4 0 0 0 0 156 0 0 503 2
640 775
229 775
2 0 5 0 0 0 0 156 0 0 504 2
640 766
166 766
1 0 6 0 0 0 0 156 0 0 505 2
640 757
99 757
2 0 167 0 0 0 0 157 0 0 486 2
635 722
514 722
5 1 168 0 0 8320 0 158 157 0 0 3
634 675
635 675
635 704
4 0 162 0 0 0 0 158 0 0 501 2
589 689
390 689
3 0 165 0 0 0 0 158 0 0 502 2
589 680
304 680
2 0 157 0 0 0 0 158 0 0 492 2
589 671
273 671
1 0 5 0 0 0 0 158 0 0 504 2
589 662
166 662
2 0 155 0 0 0 0 160 0 0 500 2
636 632
473 632
5 1 169 0 0 8320 0 159 160 0 0 4
627 584
632 584
632 614
636 614
4 0 165 0 0 0 0 159 0 0 502 2
582 598
304 598
3 0 4 0 0 0 0 159 0 0 503 2
582 589
229 589
2 0 5 0 0 0 0 159 0 0 504 2
582 580
166 580
1 0 158 0 0 0 0 159 0 0 489 2
582 571
124 571
2 0 167 0 0 0 0 162 0 0 486 2
628 532
514 532
1 0 160 0 0 0 0 162 0 0 490 2
628 514
429 514
3 0 156 0 0 0 0 163 0 0 491 2
627 488
343 488
2 0 5 0 0 0 0 163 0 0 504 2
627 479
166 479
1 0 158 0 0 0 0 163 0 0 489 2
627 470
124 470
2 3 170 0 0 8320 0 164 165 0 0 4
695 402
679 402
679 428
671 428
2 0 155 0 0 0 0 165 0 0 500 2
626 437
471 437
1 0 158 0 0 0 0 165 0 0 489 2
626 419
124 419
3 1 171 0 0 8320 0 167 166 0 0 4
624 338
615 338
615 362
623 362
2 0 162 0 0 0 0 166 0 0 501 2
623 380
390 380
2 0 165 0 0 0 0 167 0 0 502 4
575 347
309 347
309 350
304 350
1 0 4 0 0 0 0 167 0 0 503 4
575 329
245 329
245 331
230 331
3 1 172 0 0 8320 0 170 169 0 0 3
655 193
655 195
684 195
2 0 167 0 0 0 0 170 0 0 486 4
610 202
529 202
529 214
514 214
3 1 173 0 0 8320 0 177 170 0 0 3
611 181
610 181
610 184
0 2 163 0 0 0 0 0 168 493 0 4
200 281
215 281
215 237
588 237
1 0 158 0 0 0 0 168 0 0 489 4
588 219
139 219
139 263
124 263
2 0 162 0 0 0 0 177 0 0 501 2
562 190
390 190
1 0 165 0 0 0 0 177 0 0 502 2
562 172
304 172
0 2 167 0 0 8320 0 0 171 0 0 4
515 3472
514 3472
514 154
513 154
2 0 160 0 0 0 0 172 0 0 490 3
430 162
435 162
435 157
2 0 156 0 0 0 0 173 0 0 491 4
342 156
342 153
342 153
342 166
0 2 158 0 0 8320 0 0 176 0 0 3
136 3462
124 3462
124 152
0 1 160 0 0 4224 0 0 0 0 0 4
429 3470
429 162
435 162
435 154
1 0 156 0 0 12416 0 0 0 488 0 4
342 153
342 166
343 166
343 3468
2 0 157 0 0 4224 0 174 0 0 0 3
273 158
273 3468
269 3468
2 0 163 0 0 8320 0 175 0 0 0 3
199 157
200 157
200 3463
1 0 155 0 0 0 0 171 0 0 500 3
513 118
513 106
470 106
1 0 162 0 0 0 0 172 0 0 501 5
430 126
430 109
395 109
395 116
390 116
1 0 165 0 0 0 0 173 0 0 502 3
342 120
342 109
308 109
1 0 4 0 0 0 0 174 0 0 503 3
273 122
273 109
230 109
1 0 5 0 0 0 0 175 0 0 504 3
199 121
199 109
165 109
1 0 6 0 0 0 0 176 0 0 505 5
124 116
124 110
99 110
99 115
94 115
1 0 155 0 0 20608 0 7 0 0 0 6
470 101
470 151
471 151
471 437
473 437
473 3444
0 1 162 0 0 8320 0 0 8 0 0 5
389 3440
390 3440
390 112
392 112
392 104
1 0 165 0 0 12416 0 9 0 0 0 5
308 101
308 116
304 116
304 3438
305 3438
1 0 4 0 0 0 0 10 0 0 0 5
234 94
230 94
230 331
229 331
229 3438
1 0 5 0 0 0 0 11 0 0 0 5
160 97
165 97
165 148
166 148
166 3436
1 0 6 0 0 0 0 12 0 0 0 6
82 97
82 112
94 112
94 115
99 115
99 3433
56
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
2341 432 2538 456
2351 440 2527 456
22 S2'B(S0 xor Cin xor A)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
2330 273 2503 297
2340 281 2492 297
19 S2'S1'B'(Cin XOR A)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2044 158 2081 182
2054 166 2070 182
2 B'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1968 158 2005 182
1978 166 1994 182
2 A'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1877 157 1930 181
1887 165 1919 181
4 Cin'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1807 161 1852 185
1817 169 1841 185
3 S0'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1733 161 1778 185
1743 169 1767 185
3 S1'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1655 160 1700 184
1665 168 1689 184
3 S2'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1625 1396 1660 1419
1635 1406 1649 1421
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1690 1397 1729 1420
1702 1407 1716 1422
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1754 1401 1795 1424
1767 1411 1781 1426
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1824 1398 1870 1421
1836 1408 1857 1423
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1917 1400 1950 1423
1929 1410 1937 1425
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1999 1398 2034 1421
2012 1408 2020 1423
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2558 3097 2593 3120
2571 3107 2579 3122
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2476 3099 2509 3122
2488 3109 2496 3124
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2383 3097 2429 3120
2395 3107 2416 3122
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2313 3100 2354 3123
2326 3110 2340 3125
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2249 3096 2288 3119
2261 3106 2275 3121
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2184 3095 2219 3118
2194 3105 2208 3120
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2214 1859 2259 1883
2224 1867 2248 1883
3 S2'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2292 1860 2337 1884
2302 1868 2326 1884
3 S1'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2366 1860 2411 1884
2376 1868 2400 1884
3 S0'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
2436 1856 2489 1880
2446 1864 2478 1880
4 Cin'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2527 1857 2564 1881
2537 1865 2553 1881
2 A'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2603 1857 2640 1881
2613 1865 2629 1881
2 B'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
2889 1972 3062 1996
2899 1980 3051 1996
19 S2'S1'B'(Cin XOR A)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
2900 2131 3097 2155
2910 2139 3086 2155
22 S2'B(S0 xor Cin xor A)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
1346 2057 1543 2081
1356 2065 1532 2081
22 S2'B(S0 xor Cin xor A)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
1335 1898 1508 1922
1345 1906 1497 1922
19 S2'S1'B'(Cin XOR A)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1049 1783 1086 1807
1059 1791 1075 1807
2 B'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
973 1783 1010 1807
983 1791 999 1807
2 A'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
882 1782 935 1806
892 1790 924 1806
4 Cin'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
812 1786 857 1810
822 1794 846 1810
3 S0'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
738 1786 783 1810
748 1794 772 1810
3 S1'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
660 1785 705 1809
670 1793 694 1809
3 S2'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
630 3021 665 3044
640 3031 654 3046
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
695 3022 734 3045
707 3032 721 3047
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
759 3026 800 3049
772 3036 786 3051
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
829 3023 875 3046
841 3033 862 3048
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
922 3025 955 3048
934 3035 942 3050
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1004 3023 1039 3046
1017 3033 1025 3048
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
445 1324 480 1347
458 1334 466 1349
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
363 1326 396 1349
375 1336 383 1351
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
270 1324 316 1347
282 1334 303 1349
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
200 1327 241 1350
213 1337 227 1352
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
136 1323 175 1346
148 1333 162 1348
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
71 1322 106 1345
81 1332 95 1347
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
101 86 146 110
111 94 135 110
3 S2'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
179 87 224 111
189 95 213 111
3 S1'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
253 87 298 111
263 95 287 111
3 S0'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
323 83 376 107
333 91 365 107
4 Cin'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
414 84 451 108
424 92 440 108
2 A'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
490 84 527 108
500 92 516 108
2 B'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
776 199 949 223
786 207 938 223
19 S2'S1'B'(Cin XOR A)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
787 358 984 382
797 366 973 382
22 S2'B(S0 xor Cin xor A)
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
