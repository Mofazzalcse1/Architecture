CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
60 0 30 80 10
176 80 1364 699
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.499192 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
48
5 4030~
219 693 204 0 3 22
0 23 19 47
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
5130 0 0
2
44771 47
0
9 Inverter~
13 236 157 0 2 22
0 37 15
0
0 0 608 270
5 74F04
-18 -19 17 -11
3 U2A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
391 0 0
2
44771 46
0
9 Inverter~
13 311 162 0 2 22
0 14 21
0
0 0 608 270
5 74F04
-18 -19 17 -11
3 U2B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3124 0 0
2
44771 45
0
9 Inverter~
13 385 163 0 2 22
0 20 13
0
0 0 608 270
5 74F04
-18 -19 17 -11
3 U2C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
3421 0 0
2
44771 44
0
9 Inverter~
13 454 161 0 2 22
0 23 12
0
0 0 608 270
5 74F04
-18 -19 17 -11
3 U2D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
8157 0 0
2
44771 43
0
9 Inverter~
13 542 167 0 2 22
0 19 17
0
0 0 608 270
5 74F04
-18 -19 17 -11
3 U2E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
5572 0 0
2
44771 42
0
9 Inverter~
13 625 159 0 2 22
0 11 36
0
0 0 608 270
5 74F04
-18 -19 17 -11
3 U2F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
8901 0 0
2
44771 41
0
9 2-In AND~
219 767 228 0 3 22
0 47 36 46
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7361 0 0
2
44771 40
0
9 2-In AND~
219 873 257 0 3 22
0 46 45 35
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
4747 0 0
2
44771 39
0
9 2-In AND~
219 771 295 0 3 22
0 15 21 45
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
972 0 0
2
44771 38
0
5 4030~
219 692 363 0 3 22
0 20 23 44
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
3472 0 0
2
44771 37
0
5 4030~
219 754 394 0 3 22
0 44 19 43
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U1C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
9998 0 0
2
44771 36
0
9 2-In AND~
219 765 451 0 3 22
0 15 11 42
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3536 0 0
2
44771 35
0
9 2-In AND~
219 874 418 0 3 22
0 43 42 32
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
4597 0 0
2
44771 34
0
5 7415~
219 766 502 0 4 22
0 15 14 12 41
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 6 0
1 U
3835 0 0
2
44771 33
0
9 2-In AND~
219 767 546 0 3 22
0 17 36 40
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3670 0 0
2
44771 32
0
9 2-In AND~
219 879 523 0 3 22
0 41 40 33
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
5616 0 0
2
44771 31
0
9 2-In AND~
219 775 646 0 3 22
0 39 11 34
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
9323 0 0
2
44771 30
0
9 4-In AND~
219 721 607 0 5 22
0 15 14 20 23 39
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 U7A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 7 0
1 U
317 0 0
2
44771 29
0
9 4-In AND~
219 728 698 0 5 22
0 14 13 23 19 38
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 U7B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 7 0
1 U
3108 0 0
2
44771 28
0
9 2-In AND~
219 774 736 0 3 22
0 38 36 31
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
4299 0 0
2
44771 27
0
9 4-In AND~
219 779 793 0 5 22
0 37 14 20 19 28
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 U8A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 8 0
1 U
9672 0 0
2
44771 26
0
9 4-In AND~
219 781 858 0 5 22
0 37 13 17 11 30
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 U8B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 8 0
1 U
7876 0 0
2
44771 25
0
9 4-In AND~
219 781 917 0 5 22
0 49 13 19 36 29
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 U9A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 512 2 1 9 0
1 U
6369 0 0
2
44771 24
0
9 4-In AND~
219 782 977 0 5 22
0 37 21 17 48 26
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 U9B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 512 2 2 9 0
1 U
9172 0 0
2
44771 23
0
8 4-In OR~
219 991 474 0 5 22
0 35 32 33 34 25
0
0 0 608 0
4 4072
-14 -24 14 -16
4 U10A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 10 0
1 U
7100 0 0
2
44771 22
0
8 4-In OR~
219 930 793 0 5 22
0 31 28 30 29 27
0
0 0 608 0
4 4072
-14 -24 14 -16
4 U10B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 10 0
1 U
3820 0 0
2
44771 21
0
8 3-In OR~
219 1212 618 0 4 22
0 25 27 26 24
0
0 0 608 0
4 4075
-14 -24 14 -16
4 U11A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 11 0
1 U
7678 0 0
2
44771 20
0
14 Logic Display~
6 1300 603 0 1 2
10 24
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
44771 19
0
9 4-In AND~
219 780 1068 0 5 22
0 15 21 23 19 5
0
0 0 608 0
6 74LS21
-21 -28 21 -20
4 U12A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 12 0
1 U
3178 0 0
2
44771 18
0
9 4-In AND~
219 784 1142 0 5 22
0 15 21 20 23 22
0
0 0 608 0
6 74LS21
-21 -28 21 -20
4 U12B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 12 0
1 U
3409 0 0
2
44771 17
0
9 4-In AND~
219 791 1268 0 5 22
0 15 21 20 19 18
0
0 0 608 0
6 74LS21
-21 -28 21 -20
4 U13A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 13 0
1 U
3951 0 0
2
44771 16
0
9 4-In AND~
219 766 1398 0 5 22
0 15 14 12 17 8
0
0 0 608 0
6 74LS21
-21 -28 21 -20
4 U13B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 13 0
1 U
8885 0 0
2
44771 15
0
9 4-In AND~
219 790 1498 0 5 22
0 15 14 13 17 16
0
0 0 608 0
6 74LS21
-21 -28 21 -20
4 U14A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 14 0
1 U
3780 0 0
2
44771 14
0
9 4-In AND~
219 795 1610 0 5 22
0 15 14 13 12 10
0
0 0 608 0
6 74LS21
-21 -28 21 -20
4 U14B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 14 0
1 U
9265 0 0
2
44771 13
0
9 2-In AND~
219 850 1180 0 3 22
0 22 11 4
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
9442 0 0
2
44771 12
0
9 2-In AND~
219 846 1301 0 3 22
0 18 11 9
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
9424 0 0
2
44771 11
0
9 2-In AND~
219 874 1540 0 3 22
0 16 11 6
0
0 0 608 0
5 74F08
-18 -24 17 -16
4 U15A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
9968 0 0
2
44771 10
0
9 2-In AND~
219 849 1653 0 3 22
0 10 11 7
0
0 0 608 0
5 74F08
-18 -24 17 -16
4 U15B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 15 0
1 U
9281 0 0
2
44771 9
0
8 4-In OR~
219 1085 1515 0 5 22
0 9 8 6 7 3
0
0 0 608 0
4 4072
-14 -24 14 -16
4 U16A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 16 0
1 U
8464 0 0
2
44771 8
0
8 3-In OR~
219 1281 1178 0 4 22
0 5 4 3 2
0
0 0 608 0
4 4075
-14 -24 14 -16
4 U11B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 11 0
1 U
7168 0 0
2
44771 7
0
14 Logic Display~
6 1376 1161 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3171 0 0
2
44771 6
0
13 Logic Switch~
5 197 108 0 10 11
0 37 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 S2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4139 0 0
2
44771 5
0
13 Logic Switch~
5 275 108 0 1 11
0 14
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 S1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6435 0 0
2
44771 4
0
13 Logic Switch~
5 349 105 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 S0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5283 0 0
2
44771 3
0
13 Logic Switch~
5 423 112 0 1 11
0 23
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 Cin
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6874 0 0
2
44771 2
0
13 Logic Switch~
5 507 115 0 1 11
0 19
0
0 0 21344 270
2 0V
-6 -21 8 -13
1 A
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5305 0 0
2
44771 1
0
13 Logic Switch~
5 585 112 0 1 11
0 11
0
0 0 21344 270
2 0V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
34 0 0
2
44771 0
0
123
4 1 2 0 0 16 0 41 42 0 0 5
1314 1178
1364 1178
1364 1187
1376 1187
1376 1179
5 3 3 0 0 16 0 40 41 0 0 4
1118 1515
1210 1515
1210 1187
1268 1187
3 2 4 0 0 16 0 36 41 0 0 4
871 1180
1215 1180
1215 1178
1269 1178
5 1 5 0 0 16 0 30 41 0 0 4
801 1068
1215 1068
1215 1169
1268 1169
3 3 6 0 0 16 0 38 40 0 0 6
895 1540
903 1540
903 1523
1036 1523
1036 1520
1068 1520
3 4 7 0 0 16 0 39 40 0 0 4
870 1653
1055 1653
1055 1529
1068 1529
5 2 8 0 0 16 0 33 40 0 0 4
787 1398
1055 1398
1055 1511
1068 1511
3 1 9 0 0 16 0 37 40 0 0 4
867 1301
1060 1301
1060 1502
1068 1502
5 1 10 0 0 16 0 35 39 0 0 4
816 1610
820 1610
820 1644
825 1644
2 0 11 0 0 16 0 39 0 0 118 4
825 1662
593 1662
593 1663
588 1663
4 0 12 0 0 16 0 35 0 0 109 2
771 1624
458 1624
3 0 13 0 0 16 0 35 0 0 110 2
771 1615
388 1615
2 0 14 0 0 16 0 35 0 0 122 2
771 1606
281 1606
1 0 15 0 0 16 0 35 0 0 107 2
771 1597
239 1597
5 1 16 0 0 16 0 34 38 0 0 4
811 1498
842 1498
842 1531
850 1531
2 0 11 0 0 16 0 38 0 0 118 2
850 1549
588 1549
4 0 17 0 0 16 0 34 0 0 108 2
766 1512
544 1512
3 0 13 0 0 16 0 34 0 0 110 2
766 1503
388 1503
2 0 14 0 0 16 0 34 0 0 122 2
766 1494
281 1494
1 0 15 0 0 16 0 34 0 0 107 2
766 1485
239 1485
4 0 17 0 0 16 0 33 0 0 108 4
742 1412
549 1412
549 1413
544 1413
3 0 12 0 0 16 0 33 0 0 109 2
742 1403
458 1403
2 0 14 0 0 16 0 33 0 0 122 2
742 1394
281 1394
1 0 15 0 0 16 0 33 0 0 107 2
742 1385
239 1385
5 1 18 0 0 16 0 32 37 0 0 4
812 1268
816 1268
816 1292
822 1292
2 0 11 0 0 16 0 37 0 0 118 2
822 1310
588 1310
4 0 19 0 0 16 0 32 0 0 119 2
767 1282
505 1282
3 0 20 0 0 16 0 32 0 0 121 2
767 1273
344 1273
2 0 21 0 0 16 0 32 0 0 111 2
767 1264
315 1264
1 0 15 0 0 16 0 32 0 0 107 2
767 1255
239 1255
5 1 22 0 0 16 0 31 36 0 0 4
805 1142
818 1142
818 1171
826 1171
2 0 11 0 0 16 0 36 0 0 118 2
826 1189
588 1189
4 0 23 0 0 16 0 31 0 0 120 2
760 1156
419 1156
3 0 20 0 0 16 0 31 0 0 121 2
760 1147
344 1147
2 0 21 0 0 16 0 31 0 0 111 2
760 1138
315 1138
1 0 15 0 0 16 0 31 0 0 107 2
760 1129
239 1129
4 0 19 0 0 16 0 30 0 0 119 2
756 1082
505 1082
3 0 23 0 0 16 0 30 0 0 120 2
756 1073
419 1073
2 0 21 0 0 16 0 30 0 0 111 2
756 1064
315 1064
1 0 15 0 0 16 0 30 0 0 107 2
756 1055
239 1055
4 1 24 0 0 16 0 28 29 0 0 5
1245 618
1288 618
1288 629
1300 629
1300 621
5 1 25 0 0 16 0 26 28 0 0 4
1024 474
1120 474
1120 609
1199 609
5 3 26 0 0 16 0 25 28 0 0 4
803 977
1159 977
1159 627
1199 627
5 2 27 0 0 16 0 27 28 0 0 4
963 793
1120 793
1120 618
1200 618
2 5 28 0 0 16 0 27 22 0 0 3
913 789
800 789
800 793
5 4 29 0 0 16 0 24 27 0 0 4
802 917
906 917
906 807
913 807
5 3 30 0 0 16 0 23 27 0 0 4
802 858
881 858
881 798
913 798
3 1 31 0 0 16 0 21 27 0 0 4
795 736
905 736
905 780
913 780
3 2 32 0 0 16 0 14 26 0 0 4
895 418
925 418
925 470
974 470
3 3 33 0 0 16 0 17 26 0 0 4
900 523
922 523
922 479
974 479
3 4 34 0 0 16 0 18 26 0 0 4
796 646
954 646
954 488
974 488
3 1 35 0 0 16 0 9 26 0 0 4
894 257
956 257
956 461
974 461
0 0 36 0 0 16 0 0 0 0 104 2
764 992
629 992
3 0 17 0 0 16 0 25 0 0 108 2
758 982
544 982
2 0 21 0 0 16 0 25 0 0 111 2
758 973
315 973
1 0 37 0 0 16 0 25 0 0 123 2
758 964
214 964
4 0 36 0 0 16 0 24 0 0 104 2
757 931
629 931
3 0 19 0 0 16 0 24 0 0 119 2
757 922
505 922
2 0 13 0 0 16 0 24 0 0 110 2
757 913
388 913
0 0 37 0 0 16 0 0 0 0 123 2
764 905
214 905
4 0 11 0 0 16 0 23 0 0 118 2
757 872
588 872
3 0 17 0 0 16 0 23 0 0 108 2
757 863
544 863
2 0 13 0 0 16 0 23 0 0 110 2
757 854
388 854
1 0 37 0 0 16 0 23 0 0 123 2
757 845
214 845
4 0 19 0 0 16 0 22 0 0 119 2
755 807
505 807
3 0 20 0 0 16 0 22 0 0 121 2
755 798
344 798
2 0 14 0 0 16 0 22 0 0 122 2
755 789
281 789
1 0 37 0 0 16 0 22 0 0 123 2
755 780
214 780
2 0 36 0 0 16 0 21 0 0 104 2
750 745
629 745
5 1 38 0 0 16 0 20 21 0 0 3
749 698
750 698
750 727
4 0 19 0 0 16 0 20 0 0 119 2
704 712
505 712
3 0 23 0 0 16 0 20 0 0 120 2
704 703
419 703
2 0 13 0 0 16 0 20 0 0 110 2
704 694
388 694
1 0 14 0 0 16 0 20 0 0 122 2
704 685
281 685
2 0 11 0 0 16 0 18 0 0 118 2
751 655
588 655
5 1 39 0 0 16 0 19 18 0 0 4
742 607
747 607
747 637
751 637
4 0 23 0 0 16 0 19 0 0 120 2
697 621
419 621
3 0 20 0 0 16 0 19 0 0 121 2
697 612
344 612
2 0 14 0 0 16 0 19 0 0 122 2
697 603
281 603
1 0 15 0 0 16 0 19 0 0 107 2
697 594
239 594
3 2 40 0 0 16 0 16 17 0 0 4
788 546
837 546
837 532
855 532
4 1 41 0 0 16 0 15 17 0 0 4
787 502
839 502
839 514
855 514
2 0 36 0 0 16 0 16 0 0 104 2
743 555
629 555
1 0 17 0 0 16 0 16 0 0 108 2
743 537
544 537
3 0 12 0 0 16 0 15 0 0 109 2
742 511
458 511
2 0 14 0 0 16 0 15 0 0 122 2
742 502
281 502
1 0 15 0 0 16 0 15 0 0 107 2
742 493
239 493
2 3 42 0 0 16 0 14 13 0 0 4
850 427
794 427
794 451
786 451
3 1 43 0 0 16 0 12 14 0 0 4
787 394
842 394
842 409
850 409
2 0 11 0 0 16 0 13 0 0 118 2
741 460
586 460
1 0 15 0 0 16 0 13 0 0 107 2
741 442
239 442
3 1 44 0 0 16 0 11 12 0 0 4
725 363
730 363
730 385
738 385
2 0 19 0 0 16 0 12 0 0 119 2
738 403
505 403
2 0 23 0 0 16 0 11 0 0 120 4
676 372
424 372
424 373
419 373
1 0 20 0 0 16 0 11 0 0 121 2
676 354
345 354
3 2 45 0 0 16 0 10 9 0 0 4
792 295
841 295
841 266
849 266
3 1 46 0 0 16 0 8 9 0 0 4
788 228
841 228
841 248
849 248
2 0 36 0 0 16 0 8 0 0 104 2
743 237
629 237
3 1 47 0 0 16 0 1 8 0 0 4
726 204
735 204
735 219
743 219
0 2 21 0 0 16 0 0 10 111 0 2
315 304
747 304
1 0 15 0 0 16 0 10 0 0 107 2
747 286
239 286
2 0 19 0 0 16 0 1 0 0 119 2
677 213
505 213
1 0 23 0 0 16 0 1 0 0 120 2
677 195
419 195
0 2 36 0 0 16 0 0 7 0 0 4
630 3495
629 3495
629 177
628 177
2 0 17 0 0 16 0 6 0 0 108 3
545 185
550 185
550 180
2 0 12 0 0 16 0 5 0 0 109 4
457 179
457 176
457 176
457 189
0 2 15 0 0 16 0 0 2 0 0 3
251 3485
239 3485
239 175
0 1 17 0 0 16 0 0 0 0 0 4
544 3493
544 185
550 185
550 177
1 0 12 0 0 16 0 0 0 106 0 4
457 176
457 189
458 189
458 3491
2 0 13 0 0 16 0 4 0 0 0 3
388 181
388 3491
384 3491
2 0 21 0 0 16 0 3 0 0 0 3
314 180
315 180
315 3486
1 0 11 0 0 16 0 7 0 0 118 3
628 141
628 129
585 129
1 0 19 0 0 16 0 6 0 0 119 5
545 149
545 132
510 132
510 139
505 139
1 0 23 0 0 16 0 5 0 0 120 3
457 143
457 132
423 132
1 0 20 0 0 16 0 4 0 0 121 3
388 145
388 132
345 132
1 0 14 0 0 16 0 3 0 0 122 3
314 144
314 132
280 132
1 0 37 0 0 16 0 2 0 0 123 5
239 139
239 133
214 133
214 138
209 138
1 0 11 0 0 16 0 48 0 0 0 6
585 124
585 174
586 174
586 460
588 460
588 3467
0 1 19 0 0 16 0 0 47 0 0 5
504 3463
505 3463
505 135
507 135
507 127
1 0 23 0 0 16 0 46 0 0 0 5
423 124
423 139
419 139
419 3461
420 3461
1 0 20 0 0 16 0 45 0 0 0 5
349 117
345 117
345 354
344 354
344 3461
1 0 14 0 0 16 0 44 0 0 0 5
275 120
280 120
280 171
281 171
281 3459
1 0 37 0 0 16 0 43 0 0 0 6
197 120
197 135
209 135
209 138
214 138
214 3456
14
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
902 381 1099 405
912 389 1088 405
22 S2'B(S0 xor Cin xor A)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
891 222 1064 246
901 230 1053 246
19 S2'S1'B'(Cin XOR A)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
605 107 642 131
615 115 631 131
2 B'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
529 107 566 131
539 115 555 131
2 A'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
438 106 491 130
448 114 480 130
4 Cin'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
368 110 413 134
378 118 402 134
3 S0'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
294 110 339 134
304 118 328 134
3 S1'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
216 109 261 133
226 117 250 133
3 S2'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
186 1345 221 1368
196 1355 210 1370
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
251 1346 290 1369
263 1356 277 1371
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
315 1350 356 1373
328 1360 342 1375
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
385 1347 431 1370
397 1357 418 1372
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
478 1349 511 1372
490 1359 498 1374
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
560 1347 595 1370
573 1357 581 1372
1 B
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
