CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
40 1000 30 80 10
176 80 1364 699
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.499192 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
48
13 Logic Switch~
5 455 41 0 1 11
0 11
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9442 0 0
2
5.90037e-315 0
0
13 Logic Switch~
5 377 44 0 1 11
0 19
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 A
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9424 0 0
2
5.90037e-315 0
0
13 Logic Switch~
5 293 41 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 Cin
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9968 0 0
2
5.90037e-315 0
0
13 Logic Switch~
5 219 34 0 1 11
0 20
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 S0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9281 0 0
2
5.90037e-315 0
0
13 Logic Switch~
5 145 37 0 1 11
0 14
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 S1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8464 0 0
2
5.90037e-315 0
0
13 Logic Switch~
5 67 37 0 10 11
0 37 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 S2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7168 0 0
2
5.90037e-315 0
0
14 Logic Display~
6 1246 1090 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3171 0 0
2
44748.5 0
0
8 3-In OR~
219 1151 1107 0 4 22
0 5 4 3 2
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U11B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 11 0
1 U
4139 0 0
2
44748.5 0
0
8 4-In OR~
219 955 1444 0 5 22
0 9 8 6 7 3
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U16A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 16 0
1 U
6435 0 0
2
44748.5 0
0
9 2-In AND~
219 719 1582 0 3 22
0 10 11 7
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U15B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 15 0
1 U
5283 0 0
2
44748.5 0
0
9 2-In AND~
219 744 1469 0 3 22
0 16 11 6
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U15A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
6874 0 0
2
44748.5 0
0
9 2-In AND~
219 716 1230 0 3 22
0 18 11 9
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
5305 0 0
2
44748.5 0
0
9 2-In AND~
219 720 1109 0 3 22
0 22 11 4
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
34 0 0
2
44748.5 0
0
9 4-In AND~
219 665 1539 0 5 22
0 15 14 13 12 10
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U14B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 14 0
1 U
969 0 0
2
44748.5 0
0
9 4-In AND~
219 660 1427 0 5 22
0 15 14 13 17 16
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U14A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 14 0
1 U
8402 0 0
2
44748.5 0
0
9 4-In AND~
219 636 1327 0 5 22
0 15 14 12 17 8
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U13B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 13 0
1 U
3751 0 0
2
44748.5 0
0
9 4-In AND~
219 661 1197 0 5 22
0 15 21 20 19 18
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U13A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 13 0
1 U
4292 0 0
2
44748.5 0
0
9 4-In AND~
219 654 1071 0 5 22
0 15 21 20 23 22
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U12B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 12 0
1 U
6118 0 0
2
44748.5 0
0
9 4-In AND~
219 650 997 0 5 22
0 15 21 23 19 5
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U12A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 12 0
1 U
34 0 0
2
44748.5 0
0
14 Logic Display~
6 1170 532 0 1 2
10 24
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6357 0 0
2
44748.4 0
0
8 3-In OR~
219 1082 547 0 4 22
0 25 27 26 24
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U11A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 11 0
1 U
319 0 0
2
44748.4 0
0
8 4-In OR~
219 800 722 0 5 22
0 31 28 30 29 27
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U10B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 10 0
1 U
3976 0 0
2
44748.4 0
0
8 4-In OR~
219 861 403 0 5 22
0 35 32 33 34 25
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U10A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 10 0
1 U
7634 0 0
2
44748.4 0
0
9 4-In AND~
219 652 906 0 5 22
0 37 21 17 48 26
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U9B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 512 2 2 9 0
1 U
523 0 0
2
44748.4 0
0
9 4-In AND~
219 651 846 0 5 22
0 49 13 19 36 29
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U9A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 512 2 1 9 0
1 U
6748 0 0
2
44748.4 0
0
9 4-In AND~
219 651 787 0 5 22
0 37 13 17 11 30
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U8B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 8 0
1 U
6901 0 0
2
44748.4 0
0
9 4-In AND~
219 649 722 0 5 22
0 37 14 20 19 28
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U8A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 8 0
1 U
842 0 0
2
44748.4 0
0
9 2-In AND~
219 644 665 0 3 22
0 38 36 31
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3277 0 0
2
44748.4 0
0
9 4-In AND~
219 598 627 0 5 22
0 14 13 23 19 38
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U7B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 7 0
1 U
4212 0 0
2
44748.4 0
0
9 4-In AND~
219 591 536 0 5 22
0 15 14 20 23 39
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U7A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 7 0
1 U
4720 0 0
2
44748.4 0
0
9 2-In AND~
219 645 575 0 3 22
0 39 11 34
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
5551 0 0
2
44748.4 0
0
9 2-In AND~
219 749 452 0 3 22
0 41 40 33
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
6986 0 0
2
44748.4 0
0
9 2-In AND~
219 637 475 0 3 22
0 17 36 40
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
8745 0 0
2
44748.4 0
0
5 7415~
219 636 431 0 4 22
0 15 14 12 41
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 6 0
1 U
9592 0 0
2
44748.4 0
0
9 2-In AND~
219 744 347 0 3 22
0 43 42 32
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
8748 0 0
2
5.90037e-315 0
0
9 2-In AND~
219 635 380 0 3 22
0 15 11 42
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
7168 0 0
2
5.90037e-315 0
0
5 4030~
219 624 323 0 3 22
0 44 19 43
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
631 0 0
2
5.90037e-315 0
0
5 4030~
219 562 292 0 3 22
0 20 23 44
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
9466 0 0
2
5.90037e-315 0
0
9 2-In AND~
219 641 224 0 3 22
0 15 21 45
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3266 0 0
2
5.90037e-315 0
0
9 2-In AND~
219 743 186 0 3 22
0 46 45 35
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
7693 0 0
2
5.90037e-315 0
0
9 2-In AND~
219 637 157 0 3 22
0 47 36 46
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3723 0 0
2
5.90037e-315 0
0
9 Inverter~
13 495 88 0 2 22
0 11 36
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U2F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
3440 0 0
2
5.90037e-315 0
0
9 Inverter~
13 412 96 0 2 22
0 19 17
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U2E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
6263 0 0
2
5.90037e-315 0
0
9 Inverter~
13 324 90 0 2 22
0 23 12
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U2D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
4900 0 0
2
5.90037e-315 0
0
9 Inverter~
13 255 92 0 2 22
0 20 13
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U2C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
8783 0 0
2
5.90037e-315 0
0
9 Inverter~
13 181 91 0 2 22
0 14 21
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U2B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3221 0 0
2
5.90037e-315 0
0
9 Inverter~
13 106 86 0 2 22
0 37 15
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U2A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
3215 0 0
2
5.90037e-315 0
0
5 4030~
219 563 133 0 3 22
0 23 19 47
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
7903 0 0
2
5.90037e-315 0
0
123
4 1 2 0 0 4224 0 8 7 0 0 5
1184 1107
1234 1107
1234 1116
1246 1116
1246 1108
5 3 3 0 0 8320 0 9 8 0 0 4
988 1444
1080 1444
1080 1116
1138 1116
3 2 4 0 0 4224 0 13 8 0 0 4
741 1109
1085 1109
1085 1107
1139 1107
5 1 5 0 0 4224 0 19 8 0 0 4
671 997
1085 997
1085 1098
1138 1098
3 3 6 0 0 12416 0 11 9 0 0 6
765 1469
773 1469
773 1452
906 1452
906 1449
938 1449
3 4 7 0 0 4224 0 10 9 0 0 4
740 1582
925 1582
925 1458
938 1458
5 2 8 0 0 4224 0 16 9 0 0 4
657 1327
925 1327
925 1440
938 1440
3 1 9 0 0 8320 0 12 9 0 0 4
737 1230
930 1230
930 1431
938 1431
5 1 10 0 0 8320 0 14 10 0 0 4
686 1539
690 1539
690 1573
695 1573
2 0 11 0 0 4096 0 10 0 0 118 4
695 1591
463 1591
463 1592
458 1592
4 0 12 0 0 4096 0 14 0 0 109 2
641 1553
328 1553
3 0 13 0 0 4096 0 14 0 0 110 2
641 1544
258 1544
2 0 14 0 0 4096 0 14 0 0 122 2
641 1535
151 1535
1 0 15 0 0 4096 0 14 0 0 107 2
641 1526
109 1526
5 1 16 0 0 8320 0 15 11 0 0 4
681 1427
712 1427
712 1460
720 1460
2 0 11 0 0 4096 0 11 0 0 118 2
720 1478
458 1478
4 0 17 0 0 4096 0 15 0 0 108 2
636 1441
414 1441
3 0 13 0 0 0 0 15 0 0 110 2
636 1432
258 1432
2 0 14 0 0 0 0 15 0 0 122 2
636 1423
151 1423
1 0 15 0 0 0 0 15 0 0 107 2
636 1414
109 1414
4 0 17 0 0 0 0 16 0 0 108 4
612 1341
419 1341
419 1342
414 1342
3 0 12 0 0 0 0 16 0 0 109 2
612 1332
328 1332
2 0 14 0 0 0 0 16 0 0 122 2
612 1323
151 1323
1 0 15 0 0 0 0 16 0 0 107 2
612 1314
109 1314
5 1 18 0 0 8320 0 17 12 0 0 4
682 1197
686 1197
686 1221
692 1221
2 0 11 0 0 0 0 12 0 0 118 2
692 1239
458 1239
4 0 19 0 0 4096 0 17 0 0 119 2
637 1211
375 1211
3 0 20 0 0 4096 0 17 0 0 121 2
637 1202
214 1202
2 0 21 0 0 4096 0 17 0 0 111 2
637 1193
185 1193
1 0 15 0 0 0 0 17 0 0 107 2
637 1184
109 1184
5 1 22 0 0 8320 0 18 13 0 0 4
675 1071
688 1071
688 1100
696 1100
2 0 11 0 0 0 0 13 0 0 118 2
696 1118
458 1118
4 0 23 0 0 4096 0 18 0 0 120 2
630 1085
289 1085
3 0 20 0 0 0 0 18 0 0 121 2
630 1076
214 1076
2 0 21 0 0 0 0 18 0 0 111 2
630 1067
185 1067
1 0 15 0 0 0 0 18 0 0 107 2
630 1058
109 1058
4 0 19 0 0 0 0 19 0 0 119 2
626 1011
375 1011
3 0 23 0 0 0 0 19 0 0 120 2
626 1002
289 1002
2 0 21 0 0 0 0 19 0 0 111 2
626 993
185 993
1 0 15 0 0 0 0 19 0 0 107 2
626 984
109 984
4 1 24 0 0 4224 0 21 20 0 0 5
1115 547
1158 547
1158 558
1170 558
1170 550
5 1 25 0 0 8320 0 23 21 0 0 4
894 403
990 403
990 538
1069 538
5 3 26 0 0 4224 0 24 21 0 0 4
673 906
1029 906
1029 556
1069 556
5 2 27 0 0 8320 0 22 21 0 0 4
833 722
990 722
990 547
1070 547
2 5 28 0 0 4224 0 22 27 0 0 3
783 718
670 718
670 722
5 4 29 0 0 8320 0 25 22 0 0 4
672 846
776 846
776 736
783 736
5 3 30 0 0 4224 0 26 22 0 0 4
672 787
751 787
751 727
783 727
3 1 31 0 0 4224 0 28 22 0 0 4
665 665
775 665
775 709
783 709
3 2 32 0 0 8320 0 35 23 0 0 4
765 347
795 347
795 399
844 399
3 3 33 0 0 12416 0 32 23 0 0 4
770 452
792 452
792 408
844 408
3 4 34 0 0 4224 0 31 23 0 0 4
666 575
824 575
824 417
844 417
3 1 35 0 0 8320 0 40 23 0 0 4
764 186
826 186
826 390
844 390
0 0 36 0 0 4096 0 0 0 0 104 2
634 921
499 921
3 0 17 0 0 0 0 24 0 0 108 2
628 911
414 911
2 0 21 0 0 0 0 24 0 0 111 2
628 902
185 902
1 0 37 0 0 4096 0 24 0 0 123 2
628 893
84 893
4 0 36 0 0 0 0 25 0 0 104 2
627 860
499 860
3 0 19 0 0 0 0 25 0 0 119 2
627 851
375 851
2 0 13 0 0 0 0 25 0 0 110 2
627 842
258 842
0 0 37 0 0 4096 0 0 0 0 123 2
634 834
84 834
4 0 11 0 0 0 0 26 0 0 118 2
627 801
458 801
3 0 17 0 0 0 0 26 0 0 108 2
627 792
414 792
2 0 13 0 0 0 0 26 0 0 110 2
627 783
258 783
1 0 37 0 0 0 0 26 0 0 123 2
627 774
84 774
4 0 19 0 0 0 0 27 0 0 119 2
625 736
375 736
3 0 20 0 0 0 0 27 0 0 121 2
625 727
214 727
2 0 14 0 0 0 0 27 0 0 122 2
625 718
151 718
1 0 37 0 0 0 0 27 0 0 123 2
625 709
84 709
2 0 36 0 0 0 0 28 0 0 104 2
620 674
499 674
5 1 38 0 0 8320 0 29 28 0 0 3
619 627
620 627
620 656
4 0 19 0 0 0 0 29 0 0 119 2
574 641
375 641
3 0 23 0 0 0 0 29 0 0 120 2
574 632
289 632
2 0 13 0 0 0 0 29 0 0 110 2
574 623
258 623
1 0 14 0 0 0 0 29 0 0 122 2
574 614
151 614
2 0 11 0 0 0 0 31 0 0 118 2
621 584
458 584
5 1 39 0 0 8320 0 30 31 0 0 4
612 536
617 536
617 566
621 566
4 0 23 0 0 0 0 30 0 0 120 2
567 550
289 550
3 0 20 0 0 0 0 30 0 0 121 2
567 541
214 541
2 0 14 0 0 0 0 30 0 0 122 2
567 532
151 532
1 0 15 0 0 0 0 30 0 0 107 2
567 523
109 523
3 2 40 0 0 4224 0 33 32 0 0 4
658 475
707 475
707 461
725 461
4 1 41 0 0 4224 0 34 32 0 0 4
657 431
709 431
709 443
725 443
2 0 36 0 0 0 0 33 0 0 104 2
613 484
499 484
1 0 17 0 0 0 0 33 0 0 108 2
613 466
414 466
3 0 12 0 0 0 0 34 0 0 109 2
612 440
328 440
2 0 14 0 0 0 0 34 0 0 122 2
612 431
151 431
1 0 15 0 0 0 0 34 0 0 107 2
612 422
109 422
2 3 42 0 0 4224 0 35 36 0 0 4
720 356
664 356
664 380
656 380
3 1 43 0 0 4224 0 37 35 0 0 4
657 323
712 323
712 338
720 338
2 0 11 0 0 0 0 36 0 0 118 2
611 389
456 389
1 0 15 0 0 0 0 36 0 0 107 2
611 371
109 371
3 1 44 0 0 8320 0 38 37 0 0 4
595 292
600 292
600 314
608 314
2 0 19 0 0 0 0 37 0 0 119 2
608 332
375 332
2 0 23 0 0 0 0 38 0 0 120 4
546 301
294 301
294 302
289 302
1 0 20 0 0 0 0 38 0 0 121 2
546 283
215 283
3 2 45 0 0 4224 0 39 40 0 0 4
662 224
711 224
711 195
719 195
3 1 46 0 0 4224 0 41 40 0 0 4
658 157
711 157
711 177
719 177
2 0 36 0 0 0 0 41 0 0 104 2
613 166
499 166
3 1 47 0 0 8320 0 48 41 0 0 4
596 133
605 133
605 148
613 148
0 2 21 0 0 0 0 0 39 111 0 2
185 233
617 233
1 0 15 0 0 0 0 39 0 0 107 2
617 215
109 215
2 0 19 0 0 0 0 48 0 0 119 2
547 142
375 142
1 0 23 0 0 0 0 48 0 0 120 2
547 124
289 124
0 2 36 0 0 8320 0 0 42 0 0 4
500 3424
499 3424
499 106
498 106
2 0 17 0 0 0 0 43 0 0 108 3
415 114
420 114
420 109
2 0 12 0 0 0 0 44 0 0 109 4
327 108
327 105
327 105
327 118
0 2 15 0 0 8320 0 0 47 0 0 3
121 3414
109 3414
109 104
0 1 17 0 0 4224 0 0 0 0 0 4
414 3422
414 114
420 114
420 106
1 0 12 0 0 12432 0 0 0 106 0 4
327 105
327 118
328 118
328 3420
2 0 13 0 0 4224 0 45 0 0 0 3
258 110
258 3420
254 3420
2 0 21 0 0 8320 0 46 0 0 0 3
184 109
185 109
185 3415
1 0 11 0 0 0 0 42 0 0 118 3
498 70
498 58
455 58
1 0 19 0 0 0 0 43 0 0 119 5
415 78
415 61
380 61
380 68
375 68
1 0 23 0 0 0 0 44 0 0 120 3
327 72
327 61
293 61
1 0 20 0 0 0 0 45 0 0 121 3
258 74
258 61
215 61
1 0 14 0 0 0 0 46 0 0 122 3
184 73
184 61
150 61
1 0 37 0 0 0 0 47 0 0 123 5
109 68
109 62
84 62
84 67
79 67
1 0 11 0 0 20608 0 1 0 0 0 6
455 53
455 103
456 103
456 389
458 389
458 3396
0 1 19 0 0 8320 0 0 2 0 0 5
374 3392
375 3392
375 64
377 64
377 56
1 0 23 0 0 12416 0 3 0 0 0 5
293 53
293 68
289 68
289 3390
290 3390
1 0 20 0 0 16512 0 4 0 0 0 5
219 46
215 46
215 283
214 283
214 3390
1 0 14 0 0 16512 0 5 0 0 0 5
145 49
150 49
150 100
151 100
151 3388
1 0 37 0 0 20608 0 6 0 0 0 6
67 49
67 64
79 64
79 67
84 67
84 3385
14
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
430 1276 465 1299
443 1286 451 1301
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
348 1278 381 1301
360 1288 368 1303
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
255 1276 301 1299
267 1286 288 1301
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
185 1279 226 1302
198 1289 212 1304
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
121 1275 160 1298
133 1285 147 1300
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
56 1274 91 1297
66 1284 80 1299
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
86 38 131 62
96 46 120 62
3 S2'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
164 39 209 63
174 47 198 63
3 S1'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
238 39 283 63
248 47 272 63
3 S0'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
308 35 361 59
318 43 350 59
4 Cin'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
399 36 436 60
409 44 425 60
2 A'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
475 36 512 60
485 44 501 60
2 B'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
761 151 934 175
771 159 923 175
19 S2'S1'B'(Cin XOR A)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
772 310 969 334
782 318 958 334
22 S2'B(S0 xor Cin xor A)
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
