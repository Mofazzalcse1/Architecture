CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
2 80 1364 699
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.276252 0.500000
170 176 1304 347
9437202 0
0
6 Title:
5 Name:
0
0
0
65
13 Logic Switch~
5 79 81 0 1 11
0 2
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 S2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3371 0 0
2
44738.9 0
0
13 Logic Switch~
5 185 81 0 1 11
0 2
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 Cin
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7311 0 0
2
44738.9 0
0
13 Logic Switch~
5 117 81 0 1 11
0 2
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 S1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3409 0 0
2
44738.9 0
0
13 Logic Switch~
5 261 84 0 1 11
0 2
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3526 0 0
2
44738.9 0
0
13 Logic Switch~
5 217 81 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 A
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4129 0 0
2
44738.9 0
0
13 Logic Switch~
5 152 82 0 1 11
0 2
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 S0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6278 0 0
2
44738.9 0
0
14 Logic Display~
6 1267 373 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3482 0 0
2
44739 0
0
8 2-In OR~
219 1194 399 0 3 22
0 5 4 3
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U14B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 14 0
1 U
8323 0 0
2
44739 0
0
8 2-In OR~
219 1054 693 0 3 22
0 7 6 4
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U14A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
3984 0 0
2
44739 0
0
8 2-In OR~
219 839 254 0 3 22
0 13 12 5
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U13D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 13 0
1 U
7622 0 0
2
44739 0
0
8 2-In OR~
219 795 536 0 3 22
0 11 10 7
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U13C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 13 0
1 U
816 0 0
2
44739 0
0
8 2-In OR~
219 900 932 0 3 22
0 8 9 6
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U13B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
4656 0 0
2
44739 0
0
8 2-In OR~
219 541 958 0 3 22
0 19 18 15
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U13A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
6356 0 0
2
44738.9 0
0
9 2-In AND~
219 400 1108 0 3 22
0 16 17 14
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U12C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 12 0
1 U
7479 0 0
2
44738.9 0
0
9 2-In AND~
219 381 1004 0 3 22
0 21 2 20
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U12B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 12 0
1 U
5690 0 0
2
44738.9 0
0
9 2-In AND~
219 482 1032 0 3 22
0 20 2 18
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U12A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
5617 0 0
2
44738.9 0
0
9 2-In AND~
219 706 1027 0 3 22
0 15 14 9
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U10D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 10 0
1 U
3903 0 0
2
44738.9 0
0
9 2-In AND~
219 432 937 0 3 22
0 22 2 19
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U10C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
4452 0 0
2
44738.9 0
0
9 2-In AND~
219 365 895 0 3 22
0 24 23 22
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U10B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
6282 0 0
2
44738.9 0
0
9 Inverter~
13 302 911 0 2 22
0 2 23
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U11D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 11 0
1 U
7187 0 0
2
44738.9 0
0
9 Inverter~
13 309 985 0 2 22
0 2 21
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U11C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 11 0
1 U
6866 0 0
2
44738.9 0
0
9 Inverter~
13 314 1125 0 2 22
0 2 17
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U11B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 11 0
1 U
7670 0 0
2
44738.9 0
0
9 Inverter~
13 314 1095 0 2 22
0 2 16
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U11A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 11 0
1 U
951 0 0
2
44738.9 0
0
9 Inverter~
13 302 882 0 2 22
0 2 24
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U7F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 7 0
1 U
9536 0 0
2
44738.9 0
0
9 2-In AND~
219 480 781 0 3 22
0 31 2 29
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U10A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
5495 0 0
2
44738.9 0
0
9 Inverter~
13 302 843 0 2 22
0 2 27
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U7E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 7 0
1 U
8152 0 0
2
44738.9 0
0
9 Inverter~
13 302 812 0 2 22
0 2 28
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U7D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 7 0
1 U
6223 0 0
2
44738.9 0
0
9 Inverter~
13 333 732 0 2 22
0 2 32
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U7C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 7 0
1 U
5441 0 0
2
44738.9 0
0
9 Inverter~
13 300 685 0 2 22
0 2 33
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U7B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 7 0
1 U
3189 0 0
2
44738.9 0
0
9 2-In AND~
219 778 818 0 3 22
0 25 26 8
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U9D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
8460 0 0
2
44738.9 0
0
9 2-In AND~
219 423 833 0 3 22
0 28 27 26
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
5179 0 0
2
44738.9 0
0
9 2-In AND~
219 413 755 0 3 22
0 32 2 31
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
3593 0 0
2
44738.9 0
0
9 2-In AND~
219 373 694 0 3 22
0 33 2 30
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
3928 0 0
2
44738.9 0
0
8 2-In OR~
219 599 762 0 3 22
0 30 29 25
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U6D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
363 0 0
2
44738.9 0
0
8 2-In OR~
219 439 646 0 3 22
0 36 2 34
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U6C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
8132 0 0
2
44738.9 0
0
9 2-In AND~
219 333 633 0 3 22
0 2 2 36
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U8D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
65 0 0
2
44738.9 0
0
9 2-In AND~
219 560 614 0 3 22
0 35 34 10
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U8C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
6609 0 0
2
44738.9 0
0
9 2-In AND~
219 440 588 0 3 22
0 37 2 35
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U8B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
8995 0 0
2
44738.9 0
0
9 2-In AND~
219 353 551 0 3 22
0 39 38 37
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
3918 0 0
2
44738.9 0
0
9 Inverter~
13 283 563 0 2 22
0 2 38
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U7A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 7 0
1 U
7519 0 0
2
44738.9 0
0
9 Inverter~
13 283 538 0 2 22
0 2 39
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U3F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 3 0
1 U
377 0 0
2
44738.9 0
0
9 Inverter~
13 282 501 0 2 22
0 2 42
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U3E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 3 0
1 U
8816 0 0
2
44738.9 0
0
9 Inverter~
13 342 447 0 2 22
0 2 44
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U3D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
3877 0 0
2
44738.9 0
0
8 2-In OR~
219 533 449 0 3 22
0 43 2 40
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U6B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
926 0 0
2
44738.9 0
0
8 2-In OR~
219 434 436 0 3 22
0 45 44 43
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
7262 0 0
2
44738.9 0
0
9 2-In AND~
219 679 472 0 3 22
0 40 41 11
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
5267 0 0
2
44738.9 0
0
9 2-In AND~
219 396 492 0 3 22
0 2 42 41
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
8838 0 0
2
44738.9 0
0
9 2-In AND~
219 337 403 0 3 22
0 2 2 45
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
7159 0 0
2
44738.9 0
0
9 Inverter~
13 396 341 0 2 22
0 2 49
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
5812 0 0
2
44738.9 0
0
9 Inverter~
13 393 308 0 2 22
0 2 50
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
331 0 0
2
44738.9 0
0
9 2-In AND~
219 697 327 0 3 22
0 46 2 12
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
9604 0 0
2
44738.9 0
0
9 2-In AND~
219 600 300 0 3 22
0 48 47 46
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
7518 0 0
2
44738.9 0
0
9 2-In AND~
219 486 323 0 3 22
0 50 49 47
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
4832 0 0
2
44738.9 0
0
10 2-In XNOR~
219 370 276 0 3 22
0 2 2 48
0
0 0 624 0
4 4077
-7 -24 21 -16
3 U4A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
6798 0 0
2
44738.9 0
0
9 Inverter~
13 347 206 0 2 22
0 2 53
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3336 0 0
2
44738.9 0
0
9 2-In AND~
219 693 180 0 3 22
0 52 51 13
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
8370 0 0
2
44738.9 0
0
9 2-In AND~
219 548 216 0 3 22
0 53 2 51
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3910 0 0
2
44738.9 0
0
9 2-In XOR~
219 406 171 0 3 22
0 54 2 52
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
316 0 0
2
44738.9 0
0
9 2-In XOR~
219 333 126 0 3 22
0 2 2 54
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
536 0 0
2
44738.9 0
0
7 Ground~
168 249 1397 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4460 0 0
2
44738.9 0
0
7 Ground~
168 206 1397 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3260 0 0
2
44738.9 0
0
7 Ground~
168 174 1399 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5156 0 0
2
44738.9 0
0
7 Ground~
168 141 1400 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3133 0 0
2
44738.9 0
0
7 Ground~
168 111 1400 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5523 0 0
2
44738.9 0
0
7 Ground~
168 81 1402 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3746 0 0
2
44738.9 0
0
96
3 1 3 0 0 4224 0 8 7 0 0 3
1227 399
1267 399
1267 391
3 2 4 0 0 8320 0 9 8 0 0 4
1087 693
1173 693
1173 408
1181 408
3 1 5 0 0 4224 0 10 8 0 0 4
872 254
1173 254
1173 390
1181 390
3 2 6 0 0 8320 0 12 9 0 0 4
933 932
1033 932
1033 702
1041 702
3 1 7 0 0 4224 0 11 9 0 0 4
828 536
1033 536
1033 684
1041 684
3 1 8 0 0 8320 0 30 12 0 0 4
799 818
879 818
879 923
887 923
3 2 9 0 0 4224 0 17 12 0 0 4
727 1027
879 1027
879 941
887 941
3 2 10 0 0 4224 0 37 11 0 0 4
581 614
774 614
774 545
782 545
3 1 11 0 0 4224 0 46 11 0 0 4
700 472
774 472
774 527
782 527
3 2 12 0 0 4224 0 51 10 0 0 4
718 327
818 327
818 263
826 263
3 1 13 0 0 4224 0 56 10 0 0 4
714 180
818 180
818 245
826 245
3 2 14 0 0 4224 0 14 17 0 0 4
421 1108
674 1108
674 1036
682 1036
3 1 15 0 0 4224 0 13 17 0 0 4
574 958
674 958
674 1018
682 1018
2 1 16 0 0 4224 0 23 14 0 0 4
335 1095
368 1095
368 1099
376 1099
2 2 17 0 0 4224 0 22 14 0 0 4
335 1125
368 1125
368 1117
376 1117
1 0 2 0 0 4096 0 22 0 0 93 4
299 1125
179 1125
179 1126
174 1126
1 0 2 0 0 4096 0 23 0 0 96 2
299 1095
81 1095
3 2 18 0 0 8320 0 16 13 0 0 4
503 1032
520 1032
520 967
528 967
3 1 19 0 0 4224 0 18 13 0 0 4
453 937
520 937
520 949
528 949
3 1 20 0 0 4224 0 15 16 0 0 4
402 1004
450 1004
450 1023
458 1023
2 0 2 0 0 4096 0 16 0 0 95 2
458 1041
111 1041
2 1 21 0 0 4224 0 21 15 0 0 4
330 985
349 985
349 995
357 995
2 0 2 0 0 0 0 15 0 0 94 2
357 1013
141 1013
1 0 2 0 0 0 0 21 0 0 92 2
294 985
206 985
2 0 2 0 0 0 0 18 0 0 92 2
408 946
206 946
3 1 22 0 0 8320 0 19 18 0 0 4
386 895
400 895
400 928
408 928
2 2 23 0 0 4224 0 20 19 0 0 4
323 911
333 911
333 904
341 904
2 1 24 0 0 4224 0 24 19 0 0 4
323 882
333 882
333 886
341 886
1 0 2 0 0 0 0 20 0 0 94 2
287 911
141 911
1 0 2 0 0 0 0 24 0 0 95 2
287 882
111 882
3 1 25 0 0 4224 0 34 30 0 0 4
632 762
746 762
746 809
754 809
3 2 26 0 0 4224 0 31 30 0 0 4
444 833
746 833
746 827
754 827
2 2 27 0 0 4224 0 31 26 0 0 4
399 842
331 842
331 843
323 843
1 2 28 0 0 4224 0 31 27 0 0 4
399 824
331 824
331 812
323 812
1 0 2 0 0 0 0 26 0 0 91 4
287 843
254 843
254 844
249 844
1 0 2 0 0 0 0 27 0 0 95 2
287 812
111 812
3 2 29 0 0 4224 0 25 34 0 0 4
501 781
578 781
578 771
586 771
3 1 30 0 0 4224 0 33 34 0 0 4
394 694
578 694
578 753
586 753
3 1 31 0 0 8320 0 32 25 0 0 4
434 755
448 755
448 772
456 772
2 0 2 0 0 0 0 25 0 0 94 2
456 790
141 790
1 2 32 0 0 4224 0 32 28 0 0 4
389 746
362 746
362 732
354 732
2 0 2 0 0 0 0 32 0 0 92 2
389 764
206 764
1 0 2 0 0 0 0 28 0 0 44 3
318 732
271 732
271 703
2 0 2 0 0 0 0 33 0 0 93 2
349 703
174 703
1 0 2 0 0 0 0 29 0 0 92 4
285 685
211 685
211 686
206 686
2 1 33 0 0 4224 0 29 33 0 0 2
321 685
349 685
2 3 34 0 0 4224 0 37 35 0 0 4
536 623
480 623
480 646
472 646
3 1 35 0 0 4224 0 38 37 0 0 4
461 588
528 588
528 605
536 605
1 3 36 0 0 4224 0 35 36 0 0 4
426 637
362 637
362 633
354 633
2 0 2 0 0 0 0 35 0 0 96 2
426 655
81 655
2 0 2 0 0 0 0 36 0 0 93 4
309 642
179 642
179 643
174 643
1 0 2 0 0 0 0 36 0 0 95 2
309 624
111 624
2 0 2 0 0 0 0 38 0 0 92 2
416 597
206 597
3 1 37 0 0 4224 0 39 38 0 0 4
374 551
408 551
408 579
416 579
2 2 38 0 0 4224 0 39 40 0 0 4
329 560
312 560
312 563
304 563
1 2 39 0 0 4224 0 39 41 0 0 4
329 542
312 542
312 538
304 538
1 0 2 0 0 0 0 40 0 0 94 2
268 563
141 563
0 1 2 0 0 0 0 0 41 91 0 2
249 538
268 538
3 1 40 0 0 4224 0 44 46 0 0 4
566 449
647 449
647 463
655 463
3 2 41 0 0 4224 0 47 46 0 0 4
417 492
647 492
647 481
655 481
2 2 42 0 0 4224 0 47 42 0 0 2
372 501
303 501
1 0 2 0 0 0 0 42 0 0 92 2
267 501
206 501
1 0 2 0 0 0 0 47 0 0 96 2
372 483
81 483
2 0 2 0 0 0 0 44 0 0 94 4
520 458
367 458
367 462
141 462
3 1 43 0 0 4224 0 45 44 0 0 4
467 436
512 436
512 440
520 440
2 2 44 0 0 4224 0 43 45 0 0 4
363 447
413 447
413 445
421 445
0 1 2 0 0 0 0 0 43 70 0 3
284 394
284 447
327 447
3 1 45 0 0 4224 0 48 45 0 0 4
358 403
413 403
413 427
421 427
2 0 2 0 0 0 0 48 0 0 91 4
313 412
254 412
254 413
249 413
1 0 2 0 0 0 0 48 0 0 95 2
313 394
111 394
0 2 2 0 0 4096 0 0 51 95 0 4
111 358
665 358
665 336
673 336
3 1 46 0 0 4224 0 52 51 0 0 4
621 300
665 300
665 318
673 318
3 2 47 0 0 4224 0 53 52 0 0 4
507 323
568 323
568 309
576 309
1 0 48 0 0 4096 0 52 0 0 75 2
576 291
568 291
3 1 48 0 0 4224 0 54 52 0 0 4
409 276
568 276
568 291
576 291
2 2 49 0 0 4224 0 49 53 0 0 4
417 341
454 341
454 332
462 332
2 1 50 0 0 4224 0 50 53 0 0 4
414 308
454 308
454 314
462 314
1 0 2 0 0 0 0 49 0 0 96 4
381 341
86 341
86 350
81 350
1 0 2 0 0 0 0 50 0 0 92 4
378 308
221 308
221 323
206 323
2 0 2 0 0 0 0 54 0 0 91 2
354 285
249 285
1 0 2 0 0 0 0 54 0 0 93 4
354 267
179 267
179 268
174 268
3 2 51 0 0 4224 0 57 56 0 0 4
569 216
661 216
661 189
669 189
3 1 52 0 0 4224 0 58 56 0 0 2
439 171
669 171
2 0 2 0 0 0 0 57 0 0 91 2
524 225
249 225
2 1 53 0 0 4224 0 55 57 0 0 4
368 206
516 206
516 207
524 207
1 0 2 0 0 0 0 55 0 0 96 2
332 206
81 206
0 2 2 0 0 0 0 0 58 91 0 2
249 180
390 180
3 1 54 0 0 8320 0 59 58 0 0 4
366 126
382 126
382 162
390 162
0 2 2 0 0 0 0 0 59 94 0 2
141 135
317 135
1 0 2 0 0 0 0 59 0 0 93 2
317 117
174 117
1 1 2 0 0 12288 0 4 60 0 0 4
261 96
261 111
249 111
249 1391
1 1 2 0 0 12288 0 5 61 0 0 4
217 93
217 108
206 108
206 1391
1 1 2 0 0 12288 0 2 62 0 0 4
185 93
185 108
174 108
174 1393
1 1 2 0 0 0 0 6 63 0 0 4
152 94
152 109
141 109
141 1394
1 1 2 0 0 12288 0 3 64 0 0 4
117 93
117 108
111 108
111 1394
1 1 2 0 0 12416 0 1 65 0 0 4
79 93
79 108
81 108
81 1396
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1266 361 1316 376
1280 373 1301 384
3 SUM
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
